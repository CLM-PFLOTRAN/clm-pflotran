netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to patch-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to patch-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "patch-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total patch-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float RSCANOPY(time, lndgrid) ;
		RSCANOPY:long_name = "canopy resistance" ;
		RSCANOPY:units = " s m-1" ;
		RSCANOPY:cell_methods = "time: mean" ;
		RSCANOPY:_FillValue = 1.e+36f ;
		RSCANOPY:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new Patches" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total patch-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C eallocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 03/16/18 05:21:39" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "03/16/18" ;

 time_written =
  "05:21:39" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.200366e-14, 5.213594e-14, 5.211024e-14, 5.221683e-14, 5.215773e-14, 
    5.222749e-14, 5.203051e-14, 5.214117e-14, 5.207055e-14, 5.20156e-14, 
    5.242333e-14, 5.222158e-14, 5.26327e-14, 5.250429e-14, 5.282665e-14, 
    5.26127e-14, 5.286975e-14, 5.282054e-14, 5.296872e-14, 5.292629e-14, 
    5.311549e-14, 5.298829e-14, 5.321352e-14, 5.308516e-14, 5.310523e-14, 
    5.298409e-14, 5.226226e-14, 5.239821e-14, 5.225419e-14, 5.227359e-14, 
    5.226489e-14, 5.215894e-14, 5.210547e-14, 5.199357e-14, 5.20139e-14, 
    5.20961e-14, 5.228231e-14, 5.221917e-14, 5.237833e-14, 5.237474e-14, 
    5.255165e-14, 5.247192e-14, 5.276888e-14, 5.268457e-14, 5.292806e-14, 
    5.286687e-14, 5.292518e-14, 5.290751e-14, 5.292541e-14, 5.283566e-14, 
    5.287412e-14, 5.279512e-14, 5.248685e-14, 5.257752e-14, 5.230685e-14, 
    5.214371e-14, 5.203535e-14, 5.195836e-14, 5.196925e-14, 5.198999e-14, 
    5.209659e-14, 5.219676e-14, 5.227303e-14, 5.232401e-14, 5.237423e-14, 
    5.252597e-14, 5.260631e-14, 5.27859e-14, 5.275355e-14, 5.280837e-14, 
    5.286079e-14, 5.294866e-14, 5.293421e-14, 5.29729e-14, 5.280696e-14, 
    5.291726e-14, 5.273511e-14, 5.278495e-14, 5.238771e-14, 5.223621e-14, 
    5.217162e-14, 5.211518e-14, 5.197762e-14, 5.207262e-14, 5.203518e-14, 
    5.212428e-14, 5.218083e-14, 5.215287e-14, 5.23254e-14, 5.225835e-14, 
    5.261107e-14, 5.245927e-14, 5.285467e-14, 5.276019e-14, 5.287731e-14, 
    5.281757e-14, 5.29199e-14, 5.282781e-14, 5.298731e-14, 5.302199e-14, 
    5.299829e-14, 5.308936e-14, 5.28227e-14, 5.292517e-14, 5.215208e-14, 
    5.215664e-14, 5.21779e-14, 5.208441e-14, 5.20787e-14, 5.199301e-14, 
    5.206928e-14, 5.210173e-14, 5.218412e-14, 5.223281e-14, 5.227908e-14, 
    5.238074e-14, 5.249416e-14, 5.26526e-14, 5.276632e-14, 5.284247e-14, 
    5.279579e-14, 5.2837e-14, 5.279093e-14, 5.276933e-14, 5.300898e-14, 
    5.287447e-14, 5.307626e-14, 5.306511e-14, 5.297381e-14, 5.306637e-14, 
    5.215985e-14, 5.21336e-14, 5.204237e-14, 5.211377e-14, 5.198367e-14, 
    5.205649e-14, 5.209833e-14, 5.225972e-14, 5.229518e-14, 5.232801e-14, 
    5.239286e-14, 5.2476e-14, 5.26217e-14, 5.274834e-14, 5.286384e-14, 
    5.285538e-14, 5.285836e-14, 5.288413e-14, 5.282026e-14, 5.289461e-14, 
    5.290707e-14, 5.287447e-14, 5.306362e-14, 5.300962e-14, 5.306488e-14, 
    5.302972e-14, 5.214213e-14, 5.21863e-14, 5.216243e-14, 5.22073e-14, 
    5.217568e-14, 5.231617e-14, 5.235826e-14, 5.255503e-14, 5.247436e-14, 
    5.260277e-14, 5.248742e-14, 5.250786e-14, 5.260689e-14, 5.249367e-14, 
    5.274133e-14, 5.257342e-14, 5.288513e-14, 5.271761e-14, 5.289562e-14, 
    5.286334e-14, 5.291679e-14, 5.296462e-14, 5.302479e-14, 5.313568e-14, 
    5.311002e-14, 5.320272e-14, 5.225213e-14, 5.230934e-14, 5.230434e-14, 
    5.23642e-14, 5.240845e-14, 5.250434e-14, 5.265792e-14, 5.26002e-14, 
    5.270618e-14, 5.272743e-14, 5.256644e-14, 5.266528e-14, 5.234764e-14, 
    5.239899e-14, 5.236844e-14, 5.225662e-14, 5.261347e-14, 5.243046e-14, 
    5.276819e-14, 5.266923e-14, 5.29578e-14, 5.281435e-14, 5.309589e-14, 
    5.321593e-14, 5.332893e-14, 5.346066e-14, 5.234059e-14, 5.230172e-14, 
    5.237133e-14, 5.246751e-14, 5.255676e-14, 5.267526e-14, 5.26874e-14, 
    5.270957e-14, 5.276703e-14, 5.281529e-14, 5.271655e-14, 5.282739e-14, 
    5.241083e-14, 5.262935e-14, 5.2287e-14, 5.239016e-14, 5.246186e-14, 
    5.243044e-14, 5.259361e-14, 5.263203e-14, 5.278797e-14, 5.27074e-14, 
    5.318629e-14, 5.297468e-14, 5.356095e-14, 5.339743e-14, 5.228813e-14, 
    5.234047e-14, 5.252239e-14, 5.243587e-14, 5.268319e-14, 5.274396e-14, 
    5.279337e-14, 5.285645e-14, 5.286328e-14, 5.290064e-14, 5.283941e-14, 
    5.289823e-14, 5.267552e-14, 5.27751e-14, 5.250164e-14, 5.256825e-14, 
    5.253762e-14, 5.250399e-14, 5.260774e-14, 5.27181e-14, 5.272051e-14, 
    5.275586e-14, 5.285534e-14, 5.268419e-14, 5.321348e-14, 5.288683e-14, 
    5.239751e-14, 5.249813e-14, 5.251255e-14, 5.247358e-14, 5.273787e-14, 
    5.264218e-14, 5.289974e-14, 5.28302e-14, 5.294412e-14, 5.288752e-14, 
    5.287919e-14, 5.280646e-14, 5.276113e-14, 5.264656e-14, 5.255325e-14, 
    5.247924e-14, 5.249646e-14, 5.257775e-14, 5.272486e-14, 5.286388e-14, 
    5.283343e-14, 5.293547e-14, 5.266527e-14, 5.277863e-14, 5.273481e-14, 
    5.284903e-14, 5.259866e-14, 5.281175e-14, 5.254411e-14, 5.256761e-14, 
    5.264028e-14, 5.278628e-14, 5.281863e-14, 5.285307e-14, 5.283183e-14, 
    5.27286e-14, 5.27117e-14, 5.263852e-14, 5.261829e-14, 5.25625e-14, 
    5.251627e-14, 5.25585e-14, 5.260282e-14, 5.272866e-14, 5.284193e-14, 
    5.296529e-14, 5.299548e-14, 5.313928e-14, 5.302217e-14, 5.321529e-14, 
    5.305102e-14, 5.333526e-14, 5.282416e-14, 5.304629e-14, 5.26436e-14, 
    5.268707e-14, 5.276559e-14, 5.294557e-14, 5.284849e-14, 5.296204e-14, 
    5.271104e-14, 5.258053e-14, 5.25468e-14, 5.248373e-14, 5.254824e-14, 
    5.2543e-14, 5.260468e-14, 5.258487e-14, 5.273284e-14, 5.265338e-14, 
    5.287897e-14, 5.296116e-14, 5.319299e-14, 5.333483e-14, 5.347909e-14, 
    5.354268e-14, 5.356204e-14, 5.357012e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.438759e-15, -7.432297e-15, -7.433554e-15, -7.428343e-15, -7.431234e-15, 
    -7.427822e-15, -7.437451e-15, -7.432038e-15, -7.435493e-15, -7.43818e-15, 
    -7.418241e-15, -7.42811e-15, -7.408135e-15, -7.414307e-15, -7.398673e-15, 
    -7.409107e-15, -7.396572e-15, -7.398978e-15, -7.391754e-15, 
    -7.393823e-15, -7.384585e-15, -7.3908e-15, -7.379813e-15, -7.386071e-15, 
    -7.38509e-15, -7.391004e-15, -7.426128e-15, -7.419467e-15, -7.426521e-15, 
    -7.425571e-15, -7.425998e-15, -7.431173e-15, -7.433779e-15, 
    -7.439257e-15, -7.438263e-15, -7.434241e-15, -7.425144e-15, 
    -7.428233e-15, -7.420461e-15, -7.420636e-15, -7.411996e-15, 
    -7.415889e-15, -7.401498e-15, -7.405613e-15, -7.393736e-15, 
    -7.396719e-15, -7.393875e-15, -7.394738e-15, -7.393864e-15, 
    -7.398241e-15, -7.396365e-15, -7.400219e-15, -7.415159e-15, 
    -7.410833e-15, -7.423947e-15, -7.431906e-15, -7.437212e-15, 
    -7.440978e-15, -7.440445e-15, -7.439429e-15, -7.434218e-15, 
    -7.429328e-15, -7.425603e-15, -7.423113e-15, -7.420662e-15, 
    -7.413236e-15, -7.409423e-15, -7.400664e-15, -7.402247e-15, 
    -7.399568e-15, -7.397017e-15, -7.39273e-15, -7.393436e-15, -7.391547e-15, 
    -7.399642e-15, -7.394259e-15, -7.403148e-15, -7.400715e-15, 
    -7.419978e-15, -7.427401e-15, -7.430545e-15, -7.433311e-15, 
    -7.440035e-15, -7.435389e-15, -7.437219e-15, -7.43287e-15, -7.430105e-15, 
    -7.431473e-15, -7.423045e-15, -7.426319e-15, -7.409191e-15, 
    -7.416503e-15, -7.397314e-15, -7.401923e-15, -7.39621e-15, -7.399125e-15, 
    -7.394131e-15, -7.398625e-15, -7.390846e-15, -7.389152e-15, 
    -7.390309e-15, -7.385871e-15, -7.398874e-15, -7.393874e-15, 
    -7.431511e-15, -7.431288e-15, -7.43025e-15, -7.434813e-15, -7.435093e-15, 
    -7.439284e-15, -7.435556e-15, -7.433969e-15, -7.429947e-15, 
    -7.427567e-15, -7.425306e-15, -7.420341e-15, -7.414799e-15, 
    -7.407168e-15, -7.401624e-15, -7.39791e-15, -7.400188e-15, -7.398177e-15, 
    -7.400424e-15, -7.401479e-15, -7.389785e-15, -7.396346e-15, 
    -7.386509e-15, -7.387053e-15, -7.391502e-15, -7.386992e-15, 
    -7.431131e-15, -7.432415e-15, -7.43687e-15, -7.433383e-15, -7.43974e-15, 
    -7.436178e-15, -7.434131e-15, -7.426247e-15, -7.424521e-15, 
    -7.422916e-15, -7.41975e-15, -7.41569e-15, -7.408676e-15, -7.402499e-15, 
    -7.396869e-15, -7.397281e-15, -7.397136e-15, -7.395877e-15, 
    -7.398993e-15, -7.395366e-15, -7.394756e-15, -7.396348e-15, 
    -7.387126e-15, -7.389759e-15, -7.387065e-15, -7.388779e-15, 
    -7.431998e-15, -7.429839e-15, -7.431006e-15, -7.428811e-15, 
    -7.430356e-15, -7.423488e-15, -7.421432e-15, -7.411825e-15, 
    -7.415769e-15, -7.409599e-15, -7.415133e-15, -7.414133e-15, 
    -7.409388e-15, -7.414829e-15, -7.402836e-15, -7.411025e-15, 
    -7.395828e-15, -7.403987e-15, -7.395318e-15, -7.396893e-15, 
    -7.394286e-15, -7.391951e-15, -7.389019e-15, -7.383608e-15, 
    -7.384861e-15, -7.380343e-15, -7.426623e-15, -7.423825e-15, 
    -7.424074e-15, -7.42115e-15, -7.418987e-15, -7.414307e-15, -7.406911e-15, 
    -7.40973e-15, -7.40456e-15, -7.403521e-15, -7.411379e-15, -7.406549e-15, 
    -7.421955e-15, -7.419443e-15, -7.420941e-15, -7.426401e-15, 
    -7.409076e-15, -7.417907e-15, -7.401531e-15, -7.40636e-15, -7.392284e-15, 
    -7.399275e-15, -7.38555e-15, -7.379688e-15, -7.374193e-15, -7.367764e-15, 
    -7.422302e-15, -7.424202e-15, -7.420803e-15, -7.416098e-15, 
    -7.411848e-15, -7.406065e-15, -7.405475e-15, -7.404392e-15, 
    -7.401592e-15, -7.399236e-15, -7.404046e-15, -7.398646e-15, 
    -7.418854e-15, -7.408303e-15, -7.424918e-15, -7.419873e-15, 
    -7.416377e-15, -7.417913e-15, -7.410053e-15, -7.408177e-15, 
    -7.400564e-15, -7.4045e-15, -7.381131e-15, -7.391453e-15, -7.362887e-15, 
    -7.370849e-15, -7.424866e-15, -7.42231e-15, -7.413422e-15, -7.417649e-15, 
    -7.405681e-15, -7.402714e-15, -7.400306e-15, -7.397225e-15, 
    -7.396895e-15, -7.395071e-15, -7.39806e-15, -7.395191e-15, -7.406053e-15, 
    -7.401196e-15, -7.41444e-15, -7.411288e-15, -7.412684e-15, -7.414325e-15, 
    -7.409363e-15, -7.40397e-15, -7.40386e-15, -7.402131e-15, -7.397254e-15, 
    -7.405632e-15, -7.379791e-15, -7.395722e-15, -7.419524e-15, 
    -7.414602e-15, -7.413905e-15, -7.41581e-15, -7.403011e-15, -7.40768e-15, 
    -7.395116e-15, -7.398509e-15, -7.392953e-15, -7.395712e-15, 
    -7.396119e-15, -7.399667e-15, -7.401877e-15, -7.407465e-15, 
    -7.411917e-15, -7.415535e-15, -7.414693e-15, -7.410823e-15, 
    -7.403641e-15, -7.396863e-15, -7.398346e-15, -7.393375e-15, 
    -7.406554e-15, -7.401021e-15, -7.403157e-15, -7.397589e-15, 
    -7.409804e-15, -7.399385e-15, -7.412368e-15, -7.411321e-15, 
    -7.407773e-15, -7.400642e-15, -7.399073e-15, -7.39739e-15, -7.39843e-15, 
    -7.40346e-15, -7.404288e-15, -7.40786e-15, -7.408845e-15, -7.411571e-15, 
    -7.413727e-15, -7.411765e-15, -7.409599e-15, -7.40346e-15, -7.397933e-15, 
    -7.391918e-15, -7.390448e-15, -7.38342e-15, -7.389133e-15, -7.379702e-15, 
    -7.387709e-15, -7.373864e-15, -7.39879e-15, -7.387954e-15, -7.407613e-15, 
    -7.405492e-15, -7.401653e-15, -7.392872e-15, -7.397616e-15, 
    -7.392071e-15, -7.40432e-15, -7.410683e-15, -7.412235e-15, -7.415314e-15, 
    -7.412165e-15, -7.412422e-15, -7.409513e-15, -7.41048e-15, -7.403257e-15, 
    -7.407135e-15, -7.396127e-15, -7.392116e-15, -7.380815e-15, 
    -7.373898e-15, -7.366878e-15, -7.36378e-15, -7.362838e-15, -7.362444e-15 ;

 CH4_SURF_DIFF_UNSAT =
  4.975567e-14, 4.92389e-14, 4.933951e-14, 4.892169e-14, 4.915363e-14, 
    4.887982e-14, 4.965108e-14, 4.921831e-14, 4.949474e-14, 4.970927e-14, 
    4.810762e-14, 4.890303e-14, 4.72775e-14, 4.778791e-14, 4.650315e-14, 
    4.735694e-14, 4.63305e-14, 4.652794e-14, 4.593323e-14, 4.610382e-14, 
    4.534075e-14, 4.585445e-14, 4.494404e-14, 4.546361e-14, 4.53824e-14, 
    4.587135e-14, 4.874336e-14, 4.820683e-14, 4.877507e-14, 4.86987e-14, 
    4.873299e-14, 4.914881e-14, 4.935789e-14, 4.979516e-14, 4.971588e-14, 
    4.939471e-14, 4.866434e-14, 4.89127e-14, 4.828621e-14, 4.830039e-14, 
    4.760008e-14, 4.79162e-14, 4.673461e-14, 4.707126e-14, 4.609671e-14, 
    4.63423e-14, 4.610824e-14, 4.617926e-14, 4.610731e-14, 4.646737e-14, 
    4.631319e-14, 4.662971e-14, 4.785703e-14, 4.749711e-14, 4.856785e-14, 
    4.920806e-14, 4.963211e-14, 4.993225e-14, 4.988985e-14, 4.980898e-14, 
    4.939283e-14, 4.900065e-14, 4.87011e-14, 4.850041e-14, 4.830243e-14, 
    4.770145e-14, 4.738251e-14, 4.666641e-14, 4.679595e-14, 4.657651e-14, 
    4.636672e-14, 4.601382e-14, 4.607197e-14, 4.59163e-14, 4.658236e-14, 
    4.613995e-14, 4.686967e-14, 4.667038e-14, 4.824824e-14, 4.884575e-14, 
    4.909878e-14, 4.932016e-14, 4.985724e-14, 4.948653e-14, 4.963276e-14, 
    4.92847e-14, 4.90631e-14, 4.917275e-14, 4.849492e-14, 4.875877e-14, 
    4.73636e-14, 4.79661e-14, 4.63912e-14, 4.676937e-14, 4.630045e-14, 
    4.653991e-14, 4.612938e-14, 4.649889e-14, 4.585835e-14, 4.571853e-14, 
    4.581408e-14, 4.544683e-14, 4.651935e-14, 4.61082e-14, 4.917581e-14, 
    4.915793e-14, 4.907464e-14, 4.944043e-14, 4.94628e-14, 4.979732e-14, 
    4.949973e-14, 4.937279e-14, 4.905027e-14, 4.885912e-14, 4.867723e-14, 
    4.827659e-14, 4.782793e-14, 4.719843e-14, 4.674488e-14, 4.644017e-14, 
    4.66271e-14, 4.646208e-14, 4.664653e-14, 4.673293e-14, 4.577091e-14, 
    4.631173e-14, 4.54997e-14, 4.554474e-14, 4.591258e-14, 4.553967e-14, 
    4.914537e-14, 4.924824e-14, 4.960476e-14, 4.932582e-14, 4.983371e-14, 
    4.954958e-14, 4.938595e-14, 4.875319e-14, 4.861391e-14, 4.848455e-14, 
    4.822884e-14, 4.790004e-14, 4.732147e-14, 4.681664e-14, 4.635452e-14, 
    4.638843e-14, 4.637649e-14, 4.627306e-14, 4.652909e-14, 4.6231e-14, 
    4.618089e-14, 4.631183e-14, 4.555078e-14, 4.576854e-14, 4.55457e-14, 
    4.568754e-14, 4.921482e-14, 4.904168e-14, 4.913525e-14, 4.895922e-14, 
    4.908323e-14, 4.853099e-14, 4.836505e-14, 4.758642e-14, 4.79065e-14, 
    4.739672e-14, 4.785483e-14, 4.777376e-14, 4.737993e-14, 4.783013e-14, 
    4.684445e-14, 4.751311e-14, 4.626905e-14, 4.693891e-14, 4.622697e-14, 
    4.635652e-14, 4.614201e-14, 4.594963e-14, 4.570737e-14, 4.525938e-14, 
    4.536324e-14, 4.4988e-14, 4.878324e-14, 4.8558e-14, 4.85779e-14, 
    4.834192e-14, 4.816716e-14, 4.778782e-14, 4.717735e-14, 4.740713e-14, 
    4.698511e-14, 4.690024e-14, 4.754133e-14, 4.714794e-14, 4.840712e-14, 
    4.82043e-14, 4.832513e-14, 4.876545e-14, 4.735412e-14, 4.807998e-14, 
    4.673736e-14, 4.713235e-14, 4.597707e-14, 4.655252e-14, 4.542036e-14, 
    4.493399e-14, 4.447533e-14, 4.393754e-14, 4.8435e-14, 4.858819e-14, 
    4.831385e-14, 4.793341e-14, 4.757963e-14, 4.710827e-14, 4.706e-14, 
    4.69715e-14, 4.674214e-14, 4.654902e-14, 4.694346e-14, 4.650058e-14, 
    4.815711e-14, 4.729101e-14, 4.864602e-14, 4.823914e-14, 4.795589e-14, 
    4.808026e-14, 4.743338e-14, 4.728058e-14, 4.665816e-14, 4.698024e-14, 
    4.50541e-14, 4.590888e-14, 4.352722e-14, 4.419588e-14, 4.864167e-14, 
    4.843556e-14, 4.77161e-14, 4.805882e-14, 4.707679e-14, 4.683419e-14, 
    4.663678e-14, 4.638399e-14, 4.635672e-14, 4.620676e-14, 4.645243e-14, 
    4.621649e-14, 4.710726e-14, 4.670978e-14, 4.779856e-14, 4.753405e-14, 
    4.76559e-14, 4.778923e-14, 4.737722e-14, 4.693724e-14, 4.692792e-14, 
    4.678657e-14, 4.638746e-14, 4.70728e-14, 4.49433e-14, 4.626132e-14, 
    4.82105e-14, 4.781208e-14, 4.775521e-14, 4.790969e-14, 4.685853e-14, 
    4.724009e-14, 4.621043e-14, 4.648934e-14, 4.603214e-14, 4.625947e-14, 
    4.629289e-14, 4.65844e-14, 4.676561e-14, 4.72226e-14, 4.75937e-14, 
    4.788731e-14, 4.781909e-14, 4.749624e-14, 4.691031e-14, 4.635421e-14, 
    4.647617e-14, 4.606693e-14, 4.714817e-14, 4.669556e-14, 4.687061e-14, 
    4.641383e-14, 4.741321e-14, 4.656225e-14, 4.763016e-14, 4.753667e-14, 
    4.724766e-14, 4.666476e-14, 4.653567e-14, 4.639756e-14, 4.648282e-14, 
    4.689543e-14, 4.696298e-14, 4.725471e-14, 4.733512e-14, 4.7557e-14, 
    4.77406e-14, 4.757282e-14, 4.73966e-14, 4.689529e-14, 4.64422e-14, 
    4.594688e-14, 4.582549e-14, 4.524433e-14, 4.571742e-14, 4.493591e-14, 
    4.560035e-14, 4.444871e-14, 4.651296e-14, 4.562006e-14, 4.723453e-14, 
    4.706135e-14, 4.674756e-14, 4.602591e-14, 4.641598e-14, 4.595976e-14, 
    4.696563e-14, 4.748505e-14, 4.761947e-14, 4.786946e-14, 4.761375e-14, 
    4.763457e-14, 4.738937e-14, 4.746816e-14, 4.687863e-14, 4.719555e-14, 
    4.62937e-14, 4.596339e-14, 4.502732e-14, 4.4451e-14, 4.386264e-14, 
    4.360225e-14, 4.352293e-14, 4.348975e-14 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931904e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 
    1.931903e-23, 1.931904e-23, 1.931903e-23, 1.931903e-23, 1.931904e-23, 
    1.931902e-23, 1.931903e-23, 1.9319e-23, 1.931901e-23, 1.931899e-23, 
    1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931898e-23, 1.931898e-23, 1.931897e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931902e-23, 1.931902e-23, 1.931903e-23, 1.931902e-23, 
    1.931902e-23, 1.931903e-23, 1.931903e-23, 1.931904e-23, 1.931904e-23, 
    1.931903e-23, 1.931902e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 
    1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.9319e-23, 1.931901e-23, 1.931901e-23, 1.931902e-23, 
    1.931903e-23, 1.931904e-23, 1.931904e-23, 1.931904e-23, 1.931904e-23, 
    1.931903e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 1.931902e-23, 
    1.931901e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931902e-23, 1.931903e-23, 
    1.931903e-23, 1.931903e-23, 1.931904e-23, 1.931903e-23, 1.931904e-23, 
    1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931902e-23, 1.931903e-23, 
    1.9319e-23, 1.931901e-23, 1.931899e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931898e-23, 1.931899e-23, 1.931899e-23, 1.931903e-23, 
    1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931904e-23, 
    1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.9319e-23, 1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931898e-23, 
    1.931899e-23, 1.931898e-23, 1.931898e-23, 1.931899e-23, 1.931898e-23, 
    1.931903e-23, 1.931903e-23, 1.931904e-23, 1.931903e-23, 1.931904e-23, 
    1.931904e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931898e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 
    1.931903e-23, 1.931902e-23, 1.931902e-23, 1.931901e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.931901e-23, 
    1.9319e-23, 1.931901e-23, 1.931899e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931897e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 
    1.931902e-23, 1.931902e-23, 1.931901e-23, 1.9319e-23, 1.931901e-23, 
    1.9319e-23, 1.9319e-23, 1.931901e-23, 1.9319e-23, 1.931902e-23, 
    1.931902e-23, 1.931902e-23, 1.931903e-23, 1.9319e-23, 1.931902e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931898e-23, 
    1.931897e-23, 1.931897e-23, 1.931896e-23, 1.931902e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.9319e-23, 1.931899e-23, 
    1.931902e-23, 1.9319e-23, 1.931902e-23, 1.931902e-23, 1.931901e-23, 
    1.931902e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 
    1.931897e-23, 1.931898e-23, 1.931895e-23, 1.931896e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 
    1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931901e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 
    1.9319e-23, 1.931899e-23, 1.9319e-23, 1.931897e-23, 1.931899e-23, 
    1.931902e-23, 1.931901e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 
    1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 
    1.931899e-23, 1.931901e-23, 1.931899e-23, 1.931901e-23, 1.931901e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.9319e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931898e-23, 1.931898e-23, 1.931898e-23, 1.931897e-23, 
    1.931898e-23, 1.931897e-23, 1.931899e-23, 1.931898e-23, 1.9319e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.9319e-23, 1.931901e-23, 1.931901e-23, 1.931901e-23, 1.931901e-23, 
    1.931901e-23, 1.9319e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 
    1.931899e-23, 1.931899e-23, 1.931897e-23, 1.931897e-23, 1.931896e-23, 
    1.931895e-23, 1.931895e-23, 1.931895e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975319e-24, 1.975318e-24, 1.975318e-24, 1.975317e-24, 1.975317e-24, 
    1.975317e-24, 1.975318e-24, 1.975318e-24, 1.975318e-24, 1.975319e-24, 
    1.975315e-24, 1.975317e-24, 1.975314e-24, 1.975315e-24, 1.975312e-24, 
    1.975314e-24, 1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975311e-24, 
    1.97531e-24, 1.975311e-24, 1.975309e-24, 1.97531e-24, 1.97531e-24, 
    1.975311e-24, 1.975317e-24, 1.975316e-24, 1.975317e-24, 1.975317e-24, 
    1.975317e-24, 1.975317e-24, 1.975318e-24, 1.975319e-24, 1.975319e-24, 
    1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975314e-24, 1.975315e-24, 1.975313e-24, 1.975313e-24, 1.975311e-24, 
    1.975312e-24, 1.975311e-24, 1.975312e-24, 1.975311e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975315e-24, 1.975314e-24, 1.975316e-24, 
    1.975318e-24, 1.975318e-24, 1.975319e-24, 1.975319e-24, 1.975319e-24, 
    1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975311e-24, 1.975311e-24, 1.975311e-24, 1.975312e-24, 
    1.975312e-24, 1.975313e-24, 1.975313e-24, 1.975316e-24, 1.975317e-24, 
    1.975317e-24, 1.975318e-24, 1.975319e-24, 1.975318e-24, 1.975318e-24, 
    1.975318e-24, 1.975317e-24, 1.975318e-24, 1.975316e-24, 1.975317e-24, 
    1.975314e-24, 1.975315e-24, 1.975312e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975311e-24, 
    1.975311e-24, 1.97531e-24, 1.975312e-24, 1.975311e-24, 1.975318e-24, 
    1.975317e-24, 1.975317e-24, 1.975318e-24, 1.975318e-24, 1.975319e-24, 
    1.975318e-24, 1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975317e-24, 
    1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975313e-24, 1.975313e-24, 1.975311e-24, 
    1.975312e-24, 1.97531e-24, 1.97531e-24, 1.975311e-24, 1.97531e-24, 
    1.975317e-24, 1.975318e-24, 1.975318e-24, 1.975318e-24, 1.975319e-24, 
    1.975318e-24, 1.975318e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.97531e-24, 1.975311e-24, 1.97531e-24, 
    1.975311e-24, 1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975317e-24, 
    1.975317e-24, 1.975316e-24, 1.975316e-24, 1.975314e-24, 1.975315e-24, 
    1.975314e-24, 1.975315e-24, 1.975315e-24, 1.975314e-24, 1.975315e-24, 
    1.975313e-24, 1.975314e-24, 1.975312e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975311e-24, 1.97531e-24, 
    1.97531e-24, 1.975309e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975316e-24, 1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975314e-24, 
    1.975313e-24, 1.975313e-24, 1.975314e-24, 1.975314e-24, 1.975316e-24, 
    1.975316e-24, 1.975316e-24, 1.975317e-24, 1.975314e-24, 1.975315e-24, 
    1.975313e-24, 1.975313e-24, 1.975311e-24, 1.975312e-24, 1.97531e-24, 
    1.975309e-24, 1.975308e-24, 1.975307e-24, 1.975316e-24, 1.975316e-24, 
    1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975313e-24, 1.975313e-24, 1.975312e-24, 1.975313e-24, 1.975312e-24, 
    1.975316e-24, 1.975314e-24, 1.975316e-24, 1.975316e-24, 1.975315e-24, 
    1.975315e-24, 1.975314e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975309e-24, 1.975311e-24, 1.975307e-24, 1.975308e-24, 1.975316e-24, 
    1.975316e-24, 1.975315e-24, 1.975315e-24, 1.975313e-24, 1.975313e-24, 
    1.975313e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 
    1.975312e-24, 1.975313e-24, 1.975313e-24, 1.975315e-24, 1.975314e-24, 
    1.975315e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975313e-24, 1.975312e-24, 1.975313e-24, 1.975309e-24, 1.975312e-24, 
    1.975316e-24, 1.975315e-24, 1.975315e-24, 1.975315e-24, 1.975313e-24, 
    1.975314e-24, 1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975313e-24, 1.975314e-24, 1.975314e-24, 
    1.975315e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975311e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975312e-24, 1.975314e-24, 1.975312e-24, 1.975314e-24, 1.975314e-24, 
    1.975314e-24, 1.975313e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 
    1.975313e-24, 1.975313e-24, 1.975314e-24, 1.975314e-24, 1.975314e-24, 
    1.975315e-24, 1.975314e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975311e-24, 1.975311e-24, 1.97531e-24, 1.975311e-24, 1.975309e-24, 
    1.97531e-24, 1.975308e-24, 1.975312e-24, 1.975311e-24, 1.975314e-24, 
    1.975313e-24, 1.975313e-24, 1.975311e-24, 1.975312e-24, 1.975311e-24, 
    1.975313e-24, 1.975314e-24, 1.975314e-24, 1.975315e-24, 1.975314e-24, 
    1.975314e-24, 1.975314e-24, 1.975314e-24, 1.975313e-24, 1.975314e-24, 
    1.975312e-24, 1.975311e-24, 1.975309e-24, 1.975308e-24, 1.975307e-24, 
    1.975307e-24, 1.975307e-24, 1.975307e-24 ;

 CONC_CH4_SAT =
  3.549969e-08, 3.549898e-08, 3.549913e-08, 3.549852e-08, 3.549888e-08, 
    3.549846e-08, 3.549957e-08, 3.549894e-08, 3.549935e-08, 3.549965e-08, 
    3.549722e-08, 3.549849e-08, 3.549641e-08, 3.549682e-08, 3.549512e-08, 
    3.549652e-08, 3.549483e-08, 3.54952e-08, 3.549417e-08, 3.549447e-08, 
    3.549302e-08, 3.549403e-08, 3.549231e-08, 3.549329e-08, 3.549312e-08, 
    3.549406e-08, 3.549829e-08, 3.549737e-08, 3.549833e-08, 3.54982e-08, 
    3.549827e-08, 3.549886e-08, 3.549912e-08, 3.549977e-08, 3.549966e-08, 
    3.54992e-08, 3.549815e-08, 3.549854e-08, 3.549762e-08, 3.549764e-08, 
    3.549653e-08, 3.549703e-08, 3.549555e-08, 3.549612e-08, 3.549446e-08, 
    3.549488e-08, 3.549447e-08, 3.54946e-08, 3.549447e-08, 3.549509e-08, 
    3.549482e-08, 3.549538e-08, 3.549694e-08, 3.549679e-08, 3.549802e-08, 
    3.549889e-08, 3.549953e-08, 3.549995e-08, 3.549989e-08, 3.549977e-08, 
    3.549919e-08, 3.549866e-08, 3.549824e-08, 3.549793e-08, 3.549764e-08, 
    3.549662e-08, 3.549658e-08, 3.549541e-08, 3.549566e-08, 3.549526e-08, 
    3.549492e-08, 3.54943e-08, 3.549441e-08, 3.549412e-08, 3.54953e-08, 
    3.549451e-08, 3.549579e-08, 3.549545e-08, 3.549742e-08, 3.549844e-08, 
    3.549874e-08, 3.54991e-08, 3.549984e-08, 3.549933e-08, 3.549953e-08, 
    3.549907e-08, 3.549875e-08, 3.549891e-08, 3.549793e-08, 3.549831e-08, 
    3.549655e-08, 3.549709e-08, 3.549497e-08, 3.549561e-08, 3.549481e-08, 
    3.549523e-08, 3.54945e-08, 3.549516e-08, 3.549403e-08, 3.549376e-08, 
    3.549394e-08, 3.549329e-08, 3.549519e-08, 3.549446e-08, 3.549891e-08, 
    3.549889e-08, 3.549877e-08, 3.549926e-08, 3.54993e-08, 3.549977e-08, 
    3.549936e-08, 3.549917e-08, 3.549874e-08, 3.549846e-08, 3.549819e-08, 
    3.549759e-08, 3.549687e-08, 3.54963e-08, 3.549557e-08, 3.549506e-08, 
    3.549538e-08, 3.549509e-08, 3.549541e-08, 3.549556e-08, 3.549385e-08, 
    3.549481e-08, 3.549338e-08, 3.549346e-08, 3.549411e-08, 3.549346e-08, 
    3.549887e-08, 3.549902e-08, 3.54995e-08, 3.549913e-08, 3.549982e-08, 
    3.549942e-08, 3.549917e-08, 3.549827e-08, 3.54981e-08, 3.54979e-08, 
    3.549752e-08, 3.549701e-08, 3.549651e-08, 3.549568e-08, 3.549491e-08, 
    3.549497e-08, 3.549495e-08, 3.549476e-08, 3.54952e-08, 3.549469e-08, 
    3.549459e-08, 3.549483e-08, 3.549348e-08, 3.549387e-08, 3.549347e-08, 
    3.549373e-08, 3.549897e-08, 3.549872e-08, 3.549886e-08, 3.549859e-08, 
    3.549877e-08, 3.549794e-08, 3.549768e-08, 3.549647e-08, 3.549701e-08, 
    3.549662e-08, 3.549694e-08, 3.54968e-08, 3.549654e-08, 3.549691e-08, 
    3.54957e-08, 3.549678e-08, 3.549475e-08, 3.549582e-08, 3.549468e-08, 
    3.549491e-08, 3.549454e-08, 3.549419e-08, 3.549376e-08, 3.549291e-08, 
    3.549312e-08, 3.549242e-08, 3.549835e-08, 3.5498e-08, 3.549805e-08, 
    3.54977e-08, 3.549742e-08, 3.549684e-08, 3.549628e-08, 3.549667e-08, 
    3.549598e-08, 3.549583e-08, 3.549689e-08, 3.549622e-08, 3.549777e-08, 
    3.549744e-08, 3.549766e-08, 3.549831e-08, 3.549654e-08, 3.549725e-08, 
    3.549555e-08, 3.549621e-08, 3.549424e-08, 3.549521e-08, 3.549322e-08, 
    3.549226e-08, 3.549144e-08, 3.549032e-08, 3.549783e-08, 3.549807e-08, 
    3.549766e-08, 3.549703e-08, 3.549694e-08, 3.549617e-08, 3.54961e-08, 
    3.549595e-08, 3.549558e-08, 3.549524e-08, 3.549588e-08, 3.549516e-08, 
    3.549731e-08, 3.549646e-08, 3.549814e-08, 3.549749e-08, 3.549708e-08, 
    3.549728e-08, 3.549672e-08, 3.549647e-08, 3.54954e-08, 3.549598e-08, 
    3.549247e-08, 3.549408e-08, 3.548953e-08, 3.549085e-08, 3.549815e-08, 
    3.549784e-08, 3.54967e-08, 3.549725e-08, 3.549613e-08, 3.549572e-08, 
    3.54954e-08, 3.549494e-08, 3.549491e-08, 3.549464e-08, 3.549508e-08, 
    3.549467e-08, 3.549617e-08, 3.549551e-08, 3.549686e-08, 3.549686e-08, 
    3.549664e-08, 3.549685e-08, 3.549663e-08, 3.549586e-08, 3.549588e-08, 
    3.549562e-08, 3.549481e-08, 3.549613e-08, 3.549219e-08, 3.549461e-08, 
    3.54975e-08, 3.549683e-08, 3.549678e-08, 3.549703e-08, 3.549576e-08, 
    3.549639e-08, 3.549465e-08, 3.549514e-08, 3.549435e-08, 3.549474e-08, 
    3.54948e-08, 3.54953e-08, 3.549561e-08, 3.549635e-08, 3.549652e-08, 
    3.5497e-08, 3.54969e-08, 3.54968e-08, 3.549582e-08, 3.549489e-08, 
    3.549509e-08, 3.549441e-08, 3.549625e-08, 3.549547e-08, 3.549576e-08, 
    3.549501e-08, 3.549667e-08, 3.549513e-08, 3.54966e-08, 3.549688e-08, 
    3.54964e-08, 3.549539e-08, 3.549522e-08, 3.549497e-08, 3.549513e-08, 
    3.54958e-08, 3.549593e-08, 3.549642e-08, 3.549654e-08, 3.549692e-08, 
    3.549677e-08, 3.549694e-08, 3.549663e-08, 3.549582e-08, 3.549504e-08, 
    3.549417e-08, 3.549398e-08, 3.549281e-08, 3.549371e-08, 3.549216e-08, 
    3.549339e-08, 3.549127e-08, 3.549511e-08, 3.549351e-08, 3.54964e-08, 
    3.549611e-08, 3.549554e-08, 3.549428e-08, 3.549501e-08, 3.549417e-08, 
    3.549594e-08, 3.549676e-08, 3.549658e-08, 3.549697e-08, 3.549657e-08, 
    3.54966e-08, 3.549665e-08, 3.549678e-08, 3.549579e-08, 3.549633e-08, 
    3.549479e-08, 3.549419e-08, 3.549248e-08, 3.549135e-08, 3.549023e-08, 
    3.54897e-08, 3.548954e-08, 3.548947e-08,
  6.548073e-11, 6.557504e-11, 6.555676e-11, 6.563265e-11, 6.559063e-11, 
    6.564025e-11, 6.549994e-11, 6.557871e-11, 6.552849e-11, 6.548934e-11, 
    6.577938e-11, 6.563605e-11, 6.592923e-11, 6.583742e-11, 6.606719e-11, 
    6.591493e-11, 6.609787e-11, 6.6063e-11, 6.616837e-11, 6.613821e-11, 
    6.627237e-11, 6.618228e-11, 6.634209e-11, 6.625097e-11, 6.626517e-11, 
    6.617928e-11, 6.566511e-11, 6.576149e-11, 6.565935e-11, 6.567311e-11, 
    6.566698e-11, 6.559144e-11, 6.555321e-11, 6.547363e-11, 6.548812e-11, 
    6.554663e-11, 6.56793e-11, 6.563443e-11, 6.574783e-11, 6.574528e-11, 
    6.587114e-11, 6.581442e-11, 6.602626e-11, 6.596634e-11, 6.613948e-11, 
    6.609596e-11, 6.61374e-11, 6.612486e-11, 6.613757e-11, 6.607373e-11, 
    6.610108e-11, 6.604494e-11, 6.582501e-11, 6.589007e-11, 6.569683e-11, 
    6.558037e-11, 6.550337e-11, 6.544851e-11, 6.545627e-11, 6.547102e-11, 
    6.554697e-11, 6.561846e-11, 6.567282e-11, 6.570913e-11, 6.57449e-11, 
    6.585257e-11, 6.591045e-11, 6.603827e-11, 6.601539e-11, 6.605428e-11, 
    6.609163e-11, 6.615408e-11, 6.614383e-11, 6.617128e-11, 6.605337e-11, 
    6.61317e-11, 6.600231e-11, 6.603771e-11, 6.575399e-11, 6.564656e-11, 
    6.56003e-11, 6.556025e-11, 6.546222e-11, 6.55299e-11, 6.550321e-11, 
    6.556682e-11, 6.56071e-11, 6.558721e-11, 6.571012e-11, 6.566234e-11, 
    6.591385e-11, 6.580534e-11, 6.608728e-11, 6.60201e-11, 6.610339e-11, 
    6.606093e-11, 6.613361e-11, 6.606821e-11, 6.618155e-11, 6.620612e-11, 
    6.618931e-11, 6.625406e-11, 6.606456e-11, 6.613734e-11, 6.558662e-11, 
    6.558986e-11, 6.560504e-11, 6.55383e-11, 6.553424e-11, 6.547321e-11, 
    6.552758e-11, 6.555067e-11, 6.560949e-11, 6.564414e-11, 6.567709e-11, 
    6.57495e-11, 6.583015e-11, 6.594347e-11, 6.602445e-11, 6.607864e-11, 
    6.604546e-11, 6.607475e-11, 6.604198e-11, 6.602665e-11, 6.619687e-11, 
    6.61013e-11, 6.624475e-11, 6.623684e-11, 6.617191e-11, 6.623774e-11, 
    6.559215e-11, 6.557347e-11, 6.550838e-11, 6.555933e-11, 6.546656e-11, 
    6.551842e-11, 6.554818e-11, 6.56632e-11, 6.568859e-11, 6.571194e-11, 
    6.575815e-11, 6.581732e-11, 6.59215e-11, 6.601161e-11, 6.609383e-11, 
    6.608782e-11, 6.608993e-11, 6.610822e-11, 6.606282e-11, 6.611568e-11, 
    6.612448e-11, 6.610136e-11, 6.623578e-11, 6.619742e-11, 6.623668e-11, 
    6.621172e-11, 6.557956e-11, 6.561101e-11, 6.559401e-11, 6.562594e-11, 
    6.560339e-11, 6.570338e-11, 6.573332e-11, 6.587342e-11, 6.581612e-11, 
    6.590802e-11, 6.582546e-11, 6.583996e-11, 6.591071e-11, 6.582993e-11, 
    6.600652e-11, 6.5887e-11, 6.610893e-11, 6.598953e-11, 6.611639e-11, 
    6.609348e-11, 6.613148e-11, 6.616541e-11, 6.620819e-11, 6.628686e-11, 
    6.626868e-11, 6.63345e-11, 6.565792e-11, 6.569859e-11, 6.569512e-11, 
    6.573775e-11, 6.576922e-11, 6.583752e-11, 6.594732e-11, 6.590631e-11, 
    6.598172e-11, 6.59968e-11, 6.58823e-11, 6.595251e-11, 6.572588e-11, 
    6.576234e-11, 6.574073e-11, 6.566105e-11, 6.591559e-11, 6.578476e-11, 
    6.602577e-11, 6.595539e-11, 6.616056e-11, 6.605849e-11, 6.625864e-11, 
    6.634365e-11, 6.642412e-11, 6.651732e-11, 6.57209e-11, 6.569326e-11, 
    6.574285e-11, 6.581115e-11, 6.587535e-11, 6.595966e-11, 6.596835e-11, 
    6.598409e-11, 6.6025e-11, 6.605931e-11, 6.598895e-11, 6.606792e-11, 
    6.577055e-11, 6.592694e-11, 6.56827e-11, 6.575603e-11, 6.580718e-11, 
    6.578487e-11, 6.590165e-11, 6.592896e-11, 6.603978e-11, 6.598259e-11, 
    6.632258e-11, 6.61724e-11, 6.658858e-11, 6.647253e-11, 6.568358e-11, 
    6.572087e-11, 6.585026e-11, 6.578875e-11, 6.596535e-11, 6.600855e-11, 
    6.604374e-11, 6.60885e-11, 6.609342e-11, 6.611994e-11, 6.607646e-11, 
    6.611826e-11, 6.595984e-11, 6.603072e-11, 6.583563e-11, 6.588353e-11, 
    6.586124e-11, 6.58373e-11, 6.591169e-11, 6.599003e-11, 6.59919e-11, 
    6.601696e-11, 6.608718e-11, 6.596607e-11, 6.634156e-11, 6.610963e-11, 
    6.576148e-11, 6.583291e-11, 6.584334e-11, 6.581564e-11, 6.600421e-11, 
    6.593614e-11, 6.611932e-11, 6.606991e-11, 6.615089e-11, 6.611064e-11, 
    6.610471e-11, 6.605302e-11, 6.602077e-11, 6.593922e-11, 6.587228e-11, 
    6.581969e-11, 6.583194e-11, 6.589026e-11, 6.599486e-11, 6.609378e-11, 
    6.60721e-11, 6.614474e-11, 6.59526e-11, 6.603314e-11, 6.600196e-11, 
    6.608327e-11, 6.590517e-11, 6.605628e-11, 6.586585e-11, 6.588313e-11, 
    6.593479e-11, 6.603847e-11, 6.606168e-11, 6.608609e-11, 6.607107e-11, 
    6.599755e-11, 6.598559e-11, 6.593358e-11, 6.591912e-11, 6.58795e-11, 
    6.584604e-11, 6.587662e-11, 6.590808e-11, 6.599767e-11, 6.607816e-11, 
    6.616586e-11, 6.618738e-11, 6.628913e-11, 6.620605e-11, 6.634281e-11, 
    6.622615e-11, 6.642815e-11, 6.606531e-11, 6.622311e-11, 6.59372e-11, 
    6.596813e-11, 6.60238e-11, 6.61517e-11, 6.608289e-11, 6.616344e-11, 
    6.598513e-11, 6.589215e-11, 6.586776e-11, 6.582285e-11, 6.586878e-11, 
    6.586506e-11, 6.590952e-11, 6.589543e-11, 6.600064e-11, 6.594416e-11, 
    6.610451e-11, 6.616286e-11, 6.632753e-11, 6.642811e-11, 6.653061e-11, 
    6.65757e-11, 6.658943e-11, 6.659515e-11,
  3.352515e-14, 3.362234e-14, 3.360348e-14, 3.368179e-14, 3.363841e-14, 
    3.368964e-14, 3.354492e-14, 3.362613e-14, 3.357433e-14, 3.3534e-14, 
    3.383357e-14, 3.36853e-14, 3.398844e-14, 3.389359e-14, 3.413182e-14, 
    3.397361e-14, 3.416375e-14, 3.412742e-14, 3.423717e-14, 3.420574e-14, 
    3.434578e-14, 3.425168e-14, 3.441863e-14, 3.432339e-14, 3.433823e-14, 
    3.424855e-14, 3.371529e-14, 3.381506e-14, 3.370934e-14, 3.372358e-14, 
    3.371722e-14, 3.363925e-14, 3.359985e-14, 3.351783e-14, 3.353275e-14, 
    3.359305e-14, 3.372998e-14, 3.36836e-14, 3.380081e-14, 3.379816e-14, 
    3.392855e-14, 3.386975e-14, 3.408921e-14, 3.402692e-14, 3.420706e-14, 
    3.416173e-14, 3.42049e-14, 3.419183e-14, 3.420507e-14, 3.41386e-14, 
    3.416707e-14, 3.410863e-14, 3.388074e-14, 3.394778e-14, 3.374808e-14, 
    3.362789e-14, 3.354846e-14, 3.349198e-14, 3.349996e-14, 3.351515e-14, 
    3.35934e-14, 3.366712e-14, 3.372325e-14, 3.376078e-14, 3.379778e-14, 
    3.390936e-14, 3.396895e-14, 3.410172e-14, 3.40779e-14, 3.411837e-14, 
    3.415723e-14, 3.422228e-14, 3.421159e-14, 3.424022e-14, 3.41174e-14, 
    3.419898e-14, 3.406429e-14, 3.410111e-14, 3.380729e-14, 3.369614e-14, 
    3.364843e-14, 3.360709e-14, 3.350609e-14, 3.35758e-14, 3.354831e-14, 
    3.361384e-14, 3.36554e-14, 3.363487e-14, 3.37618e-14, 3.371243e-14, 
    3.397247e-14, 3.386037e-14, 3.415269e-14, 3.40828e-14, 3.416947e-14, 
    3.412527e-14, 3.420095e-14, 3.413284e-14, 3.425092e-14, 3.427657e-14, 
    3.425903e-14, 3.432659e-14, 3.412905e-14, 3.420485e-14, 3.363427e-14, 
    3.363761e-14, 3.365326e-14, 3.358446e-14, 3.358028e-14, 3.35174e-14, 
    3.35734e-14, 3.35972e-14, 3.365785e-14, 3.369363e-14, 3.372767e-14, 
    3.380254e-14, 3.388607e-14, 3.40032e-14, 3.408732e-14, 3.414369e-14, 
    3.410916e-14, 3.413964e-14, 3.410555e-14, 3.408959e-14, 3.426692e-14, 
    3.41673e-14, 3.431687e-14, 3.430862e-14, 3.424088e-14, 3.430955e-14, 
    3.363997e-14, 3.36207e-14, 3.355362e-14, 3.360612e-14, 3.351055e-14, 
    3.356398e-14, 3.359465e-14, 3.371334e-14, 3.373956e-14, 3.376369e-14, 
    3.381149e-14, 3.387276e-14, 3.398039e-14, 3.407398e-14, 3.415951e-14, 
    3.415325e-14, 3.415545e-14, 3.41745e-14, 3.412724e-14, 3.418227e-14, 
    3.419145e-14, 3.416735e-14, 3.430751e-14, 3.426747e-14, 3.430844e-14, 
    3.428239e-14, 3.362698e-14, 3.365943e-14, 3.364188e-14, 3.367485e-14, 
    3.365158e-14, 3.375488e-14, 3.378585e-14, 3.393093e-14, 3.387152e-14, 
    3.396639e-14, 3.388119e-14, 3.389623e-14, 3.396925e-14, 3.388582e-14, 
    3.406872e-14, 3.394462e-14, 3.417524e-14, 3.405109e-14, 3.418301e-14, 
    3.415914e-14, 3.419871e-14, 3.42341e-14, 3.427872e-14, 3.436088e-14, 
    3.434188e-14, 3.441068e-14, 3.370786e-14, 3.37499e-14, 3.37463e-14, 
    3.379038e-14, 3.382295e-14, 3.389368e-14, 3.400718e-14, 3.396459e-14, 
    3.404289e-14, 3.405857e-14, 3.393969e-14, 3.401258e-14, 3.377812e-14, 
    3.381586e-14, 3.379347e-14, 3.371112e-14, 3.397427e-14, 3.383906e-14, 
    3.40887e-14, 3.401556e-14, 3.422904e-14, 3.412276e-14, 3.433139e-14, 
    3.442031e-14, 3.450447e-14, 3.460226e-14, 3.377296e-14, 3.374438e-14, 
    3.379565e-14, 3.386639e-14, 3.39325e-14, 3.402e-14, 3.402901e-14, 
    3.404537e-14, 3.408788e-14, 3.412358e-14, 3.405044e-14, 3.413253e-14, 
    3.382441e-14, 3.398604e-14, 3.373348e-14, 3.380934e-14, 3.386227e-14, 
    3.383915e-14, 3.395975e-14, 3.398811e-14, 3.410328e-14, 3.40438e-14, 
    3.439827e-14, 3.424143e-14, 3.467706e-14, 3.455526e-14, 3.373437e-14, 
    3.377291e-14, 3.390691e-14, 3.384317e-14, 3.402589e-14, 3.407079e-14, 
    3.410737e-14, 3.415397e-14, 3.415908e-14, 3.418671e-14, 3.414143e-14, 
    3.418496e-14, 3.402018e-14, 3.409383e-14, 3.389172e-14, 3.394097e-14, 
    3.391826e-14, 3.389345e-14, 3.397017e-14, 3.405157e-14, 3.405348e-14, 
    3.407955e-14, 3.415272e-14, 3.402664e-14, 3.44182e-14, 3.417609e-14, 
    3.381493e-14, 3.388895e-14, 3.389972e-14, 3.387101e-14, 3.406628e-14, 
    3.399556e-14, 3.418606e-14, 3.413461e-14, 3.421895e-14, 3.417702e-14, 
    3.417085e-14, 3.411704e-14, 3.408349e-14, 3.399877e-14, 3.392973e-14, 
    3.38752e-14, 3.388789e-14, 3.394796e-14, 3.405659e-14, 3.415947e-14, 
    3.413691e-14, 3.421254e-14, 3.401265e-14, 3.409638e-14, 3.406396e-14, 
    3.414852e-14, 3.396343e-14, 3.412054e-14, 3.392305e-14, 3.394055e-14, 
    3.399416e-14, 3.410195e-14, 3.412604e-14, 3.415147e-14, 3.413581e-14, 
    3.405937e-14, 3.404693e-14, 3.39929e-14, 3.39779e-14, 3.393678e-14, 
    3.39025e-14, 3.39338e-14, 3.396645e-14, 3.405948e-14, 3.414322e-14, 
    3.423458e-14, 3.4257e-14, 3.436333e-14, 3.427654e-14, 3.441952e-14, 
    3.429761e-14, 3.450881e-14, 3.412989e-14, 3.429437e-14, 3.399666e-14, 
    3.402877e-14, 3.408667e-14, 3.421985e-14, 3.414813e-14, 3.423208e-14, 
    3.404645e-14, 3.394995e-14, 3.392502e-14, 3.387848e-14, 3.392609e-14, 
    3.392222e-14, 3.396793e-14, 3.39533e-14, 3.406257e-14, 3.400388e-14, 
    3.417065e-14, 3.423146e-14, 3.440341e-14, 3.450871e-14, 3.461616e-14, 
    3.466351e-14, 3.467793e-14, 3.468395e-14,
  5.202264e-18, 5.224354e-18, 5.220025e-18, 5.238011e-18, 5.228042e-18, 
    5.239815e-18, 5.206715e-18, 5.225228e-18, 5.21334e-18, 5.204253e-18, 
    5.272941e-18, 5.238818e-18, 5.30862e-18, 5.286758e-18, 5.341757e-18, 
    5.305199e-18, 5.349145e-18, 5.340734e-18, 5.366144e-18, 5.358862e-18, 
    5.391341e-18, 5.369506e-18, 5.408257e-18, 5.386141e-18, 5.389586e-18, 
    5.368781e-18, 5.245709e-18, 5.268678e-18, 5.244341e-18, 5.247616e-18, 
    5.246154e-18, 5.228237e-18, 5.219197e-18, 5.200613e-18, 5.203973e-18, 
    5.217633e-18, 5.24909e-18, 5.238424e-18, 5.26538e-18, 5.264772e-18, 
    5.294819e-18, 5.281263e-18, 5.331895e-18, 5.317499e-18, 5.359167e-18, 
    5.348672e-18, 5.358668e-18, 5.35564e-18, 5.358707e-18, 5.34332e-18, 
    5.349909e-18, 5.336387e-18, 5.283795e-18, 5.299232e-18, 5.253251e-18, 
    5.225635e-18, 5.207512e-18, 5.194794e-18, 5.196591e-18, 5.200011e-18, 
    5.217713e-18, 5.234636e-18, 5.247538e-18, 5.256169e-18, 5.264684e-18, 
    5.290404e-18, 5.30412e-18, 5.334793e-18, 5.32928e-18, 5.338641e-18, 
    5.34763e-18, 5.362694e-18, 5.360218e-18, 5.366852e-18, 5.338414e-18, 
    5.357299e-18, 5.326134e-18, 5.334648e-18, 5.266892e-18, 5.241305e-18, 
    5.230352e-18, 5.220853e-18, 5.197971e-18, 5.213675e-18, 5.207479e-18, 
    5.2224e-18, 5.231945e-18, 5.227228e-18, 5.256406e-18, 5.245051e-18, 
    5.304932e-18, 5.279102e-18, 5.346581e-18, 5.330413e-18, 5.350463e-18, 
    5.340234e-18, 5.357756e-18, 5.341986e-18, 5.369331e-18, 5.375279e-18, 
    5.371212e-18, 5.386879e-18, 5.341109e-18, 5.358657e-18, 5.227091e-18, 
    5.227859e-18, 5.231453e-18, 5.215661e-18, 5.214701e-18, 5.200516e-18, 
    5.21313e-18, 5.218585e-18, 5.232507e-18, 5.240729e-18, 5.248556e-18, 
    5.265782e-18, 5.285027e-18, 5.312025e-18, 5.33146e-18, 5.344496e-18, 
    5.336508e-18, 5.343559e-18, 5.335673e-18, 5.331983e-18, 5.373043e-18, 
    5.349964e-18, 5.384624e-18, 5.382708e-18, 5.367006e-18, 5.382925e-18, 
    5.228401e-18, 5.223975e-18, 5.208675e-18, 5.220628e-18, 5.198975e-18, 
    5.211008e-18, 5.218002e-18, 5.245265e-18, 5.251287e-18, 5.256841e-18, 
    5.267841e-18, 5.281956e-18, 5.306759e-18, 5.328378e-18, 5.348157e-18, 
    5.346709e-18, 5.347218e-18, 5.351629e-18, 5.340691e-18, 5.353426e-18, 
    5.355554e-18, 5.349974e-18, 5.382451e-18, 5.373167e-18, 5.382667e-18, 
    5.376625e-18, 5.225416e-18, 5.23287e-18, 5.22884e-18, 5.236413e-18, 
    5.231069e-18, 5.254817e-18, 5.261944e-18, 5.295374e-18, 5.281672e-18, 
    5.303528e-18, 5.283898e-18, 5.287366e-18, 5.304196e-18, 5.284964e-18, 
    5.327164e-18, 5.29851e-18, 5.3518e-18, 5.323094e-18, 5.353598e-18, 
    5.348071e-18, 5.357234e-18, 5.365433e-18, 5.375774e-18, 5.394841e-18, 
    5.390428e-18, 5.406405e-18, 5.243999e-18, 5.253671e-18, 5.252838e-18, 
    5.262981e-18, 5.270481e-18, 5.286778e-18, 5.312943e-18, 5.30311e-18, 
    5.321189e-18, 5.324814e-18, 5.297361e-18, 5.314192e-18, 5.260162e-18, 
    5.268854e-18, 5.263694e-18, 5.24475e-18, 5.305347e-18, 5.274197e-18, 
    5.331777e-18, 5.314876e-18, 5.364261e-18, 5.339659e-18, 5.387995e-18, 
    5.40865e-18, 5.428211e-18, 5.450987e-18, 5.258974e-18, 5.252397e-18, 
    5.264193e-18, 5.280493e-18, 5.295705e-18, 5.315902e-18, 5.317982e-18, 
    5.321763e-18, 5.331588e-18, 5.339843e-18, 5.322939e-18, 5.341915e-18, 
    5.27083e-18, 5.308062e-18, 5.249892e-18, 5.267352e-18, 5.279541e-18, 
    5.274213e-18, 5.301992e-18, 5.308536e-18, 5.335152e-18, 5.321399e-18, 
    5.403531e-18, 5.367136e-18, 5.468421e-18, 5.440038e-18, 5.250094e-18, 
    5.25896e-18, 5.289831e-18, 5.275138e-18, 5.317263e-18, 5.327637e-18, 
    5.336095e-18, 5.346879e-18, 5.348059e-18, 5.354455e-18, 5.343973e-18, 
    5.354049e-18, 5.315945e-18, 5.332964e-18, 5.286323e-18, 5.29766e-18, 
    5.292443e-18, 5.286723e-18, 5.304396e-18, 5.3232e-18, 5.323635e-18, 
    5.329664e-18, 5.346607e-18, 5.317434e-18, 5.408173e-18, 5.352014e-18, 
    5.268633e-18, 5.285692e-18, 5.288171e-18, 5.281552e-18, 5.326596e-18, 
    5.31026e-18, 5.354304e-18, 5.342395e-18, 5.361922e-18, 5.352212e-18, 
    5.350783e-18, 5.33833e-18, 5.330574e-18, 5.311002e-18, 5.295092e-18, 
    5.282516e-18, 5.285441e-18, 5.299274e-18, 5.324359e-18, 5.348151e-18, 
    5.342931e-18, 5.360437e-18, 5.314204e-18, 5.333556e-18, 5.326063e-18, 
    5.345615e-18, 5.302841e-18, 5.339158e-18, 5.293548e-18, 5.29756e-18, 
    5.309936e-18, 5.334847e-18, 5.340413e-18, 5.346299e-18, 5.342674e-18, 
    5.325002e-18, 5.322123e-18, 5.309643e-18, 5.306182e-18, 5.296692e-18, 
    5.28881e-18, 5.296004e-18, 5.303542e-18, 5.325023e-18, 5.34439e-18, 
    5.365544e-18, 5.370739e-18, 5.395418e-18, 5.37528e-18, 5.40848e-18, 
    5.38018e-18, 5.429236e-18, 5.341314e-18, 5.379416e-18, 5.31051e-18, 
    5.317926e-18, 5.331314e-18, 5.362136e-18, 5.345524e-18, 5.36497e-18, 
    5.322013e-18, 5.299735e-18, 5.294003e-18, 5.283274e-18, 5.294248e-18, 
    5.293357e-18, 5.303878e-18, 5.300502e-18, 5.325737e-18, 5.312178e-18, 
    5.350738e-18, 5.364825e-18, 5.404718e-18, 5.429202e-18, 5.454218e-18, 
    5.465257e-18, 5.468621e-18, 5.470026e-18,
  2.57814e-22, 2.592588e-22, 2.589753e-22, 2.601536e-22, 2.595002e-22, 
    2.602718e-22, 2.581047e-22, 2.593162e-22, 2.585378e-22, 2.579437e-22, 
    2.624463e-22, 2.602064e-22, 2.648164e-22, 2.633592e-22, 2.670297e-22, 
    2.645884e-22, 2.675238e-22, 2.669609e-22, 2.686613e-22, 2.681737e-22, 
    2.703513e-22, 2.688866e-22, 2.714867e-22, 2.700021e-22, 2.702334e-22, 
    2.68838e-22, 2.60658e-22, 2.621664e-22, 2.605684e-22, 2.607832e-22, 
    2.606872e-22, 2.595131e-22, 2.589215e-22, 2.577059e-22, 2.579254e-22, 
    2.588189e-22, 2.608799e-22, 2.601804e-22, 2.619486e-22, 2.619087e-22, 
    2.638963e-22, 2.629931e-22, 2.663701e-22, 2.654084e-22, 2.681941e-22, 
    2.674918e-22, 2.681608e-22, 2.679581e-22, 2.681634e-22, 2.671339e-22, 
    2.675746e-22, 2.666703e-22, 2.631618e-22, 2.6419e-22, 2.611528e-22, 
    2.593432e-22, 2.581568e-22, 2.573258e-22, 2.574432e-22, 2.576667e-22, 
    2.588241e-22, 2.599322e-22, 2.607778e-22, 2.613441e-22, 2.619029e-22, 
    2.636028e-22, 2.645162e-22, 2.66564e-22, 2.661953e-22, 2.668212e-22, 
    2.67422e-22, 2.684304e-22, 2.682645e-22, 2.687089e-22, 2.668058e-22, 
    2.680693e-22, 2.65985e-22, 2.66554e-22, 2.620491e-22, 2.603693e-22, 
    2.596521e-22, 2.590296e-22, 2.575333e-22, 2.585598e-22, 2.581547e-22, 
    2.591307e-22, 2.597558e-22, 2.594468e-22, 2.613596e-22, 2.606148e-22, 
    2.645704e-22, 2.628503e-22, 2.673519e-22, 2.66271e-22, 2.676116e-22, 
    2.669274e-22, 2.680998e-22, 2.670445e-22, 2.688749e-22, 2.692737e-22, 
    2.69001e-22, 2.700513e-22, 2.669859e-22, 2.681602e-22, 2.594378e-22, 
    2.594882e-22, 2.597236e-22, 2.586898e-22, 2.586269e-22, 2.576996e-22, 
    2.585241e-22, 2.588811e-22, 2.597926e-22, 2.603314e-22, 2.608447e-22, 
    2.619751e-22, 2.63244e-22, 2.650434e-22, 2.66341e-22, 2.672124e-22, 
    2.666783e-22, 2.671498e-22, 2.666225e-22, 2.663758e-22, 2.691238e-22, 
    2.675784e-22, 2.699001e-22, 2.697715e-22, 2.687193e-22, 2.69786e-22, 
    2.595237e-22, 2.592338e-22, 2.582328e-22, 2.590146e-22, 2.575989e-22, 
    2.583854e-22, 2.588431e-22, 2.606291e-22, 2.610238e-22, 2.613882e-22, 
    2.621102e-22, 2.630392e-22, 2.64692e-22, 2.661352e-22, 2.674573e-22, 
    2.673604e-22, 2.673944e-22, 2.676896e-22, 2.66958e-22, 2.678099e-22, 
    2.679524e-22, 2.675789e-22, 2.697543e-22, 2.691319e-22, 2.697688e-22, 
    2.693636e-22, 2.593281e-22, 2.598164e-22, 2.595524e-22, 2.600486e-22, 
    2.596985e-22, 2.612557e-22, 2.617236e-22, 2.639336e-22, 2.630204e-22, 
    2.644766e-22, 2.631685e-22, 2.633997e-22, 2.645217e-22, 2.632395e-22, 
    2.660544e-22, 2.641423e-22, 2.677011e-22, 2.657828e-22, 2.678214e-22, 
    2.674515e-22, 2.680647e-22, 2.686138e-22, 2.693067e-22, 2.705858e-22, 
    2.702896e-22, 2.713621e-22, 2.605458e-22, 2.611803e-22, 2.611255e-22, 
    2.617912e-22, 2.622838e-22, 2.633603e-22, 2.651045e-22, 2.644484e-22, 
    2.656548e-22, 2.65897e-22, 2.64065e-22, 2.65188e-22, 2.616063e-22, 
    2.621773e-22, 2.61838e-22, 2.605952e-22, 2.64598e-22, 2.625282e-22, 
    2.663622e-22, 2.652334e-22, 2.685353e-22, 2.668893e-22, 2.701263e-22, 
    2.715135e-22, 2.728279e-22, 2.74362e-22, 2.615282e-22, 2.610965e-22, 
    2.618707e-22, 2.629422e-22, 2.639548e-22, 2.65302e-22, 2.654407e-22, 
    2.656932e-22, 2.663494e-22, 2.669012e-22, 2.65772e-22, 2.670397e-22, 
    2.623076e-22, 2.64779e-22, 2.609324e-22, 2.620787e-22, 2.628791e-22, 
    2.625289e-22, 2.643737e-22, 2.648103e-22, 2.665879e-22, 2.656688e-22, 
    2.711698e-22, 2.687283e-22, 2.755369e-22, 2.736243e-22, 2.609455e-22, 
    2.615272e-22, 2.63564e-22, 2.625896e-22, 2.653927e-22, 2.660856e-22, 
    2.666506e-22, 2.67372e-22, 2.674507e-22, 2.678789e-22, 2.671774e-22, 
    2.678515e-22, 2.653049e-22, 2.664415e-22, 2.6333e-22, 2.640851e-22, 
    2.637377e-22, 2.633566e-22, 2.645341e-22, 2.657895e-22, 2.658182e-22, 
    2.662211e-22, 2.673552e-22, 2.654041e-22, 2.714824e-22, 2.677167e-22, 
    2.621622e-22, 2.632885e-22, 2.634532e-22, 2.630122e-22, 2.66016e-22, 
    2.649254e-22, 2.678687e-22, 2.670719e-22, 2.683786e-22, 2.677286e-22, 
    2.67633e-22, 2.668001e-22, 2.662818e-22, 2.64975e-22, 2.639145e-22, 
    2.630764e-22, 2.632712e-22, 2.641928e-22, 2.658668e-22, 2.674571e-22, 
    2.67108e-22, 2.682792e-22, 2.651885e-22, 2.664812e-22, 2.659806e-22, 
    2.672873e-22, 2.644306e-22, 2.668568e-22, 2.638113e-22, 2.640783e-22, 
    2.649038e-22, 2.665678e-22, 2.669394e-22, 2.673332e-22, 2.670905e-22, 
    2.659097e-22, 2.657173e-22, 2.648841e-22, 2.646534e-22, 2.640204e-22, 
    2.634957e-22, 2.639746e-22, 2.644774e-22, 2.65911e-22, 2.672055e-22, 
    2.686214e-22, 2.689692e-22, 2.706253e-22, 2.692743e-22, 2.715031e-22, 
    2.696039e-22, 2.72898e-22, 2.670004e-22, 2.695517e-22, 2.64942e-22, 
    2.65437e-22, 2.663316e-22, 2.683935e-22, 2.672812e-22, 2.685832e-22, 
    2.657099e-22, 2.642237e-22, 2.638417e-22, 2.631269e-22, 2.638581e-22, 
    2.637986e-22, 2.644995e-22, 2.642744e-22, 2.659587e-22, 2.650533e-22, 
    2.676301e-22, 2.685734e-22, 2.71249e-22, 2.728951e-22, 2.745791e-22, 
    2.753233e-22, 2.755502e-22, 2.75645e-22,
  4.167635e-27, 4.196607e-27, 4.190941e-27, 4.214522e-27, 4.201429e-27, 
    4.216913e-27, 4.173481e-27, 4.197756e-27, 4.182198e-27, 4.170241e-27, 
    4.260971e-27, 4.215589e-27, 4.309129e-27, 4.279485e-27, 4.354246e-27, 
    4.304491e-27, 4.36433e-27, 4.352834e-27, 4.387567e-27, 4.377599e-27, 
    4.422168e-27, 4.392173e-27, 4.445438e-27, 4.415008e-27, 4.419748e-27, 
    4.391181e-27, 4.224722e-27, 4.255295e-27, 4.222909e-27, 4.22726e-27, 
    4.225313e-27, 4.201689e-27, 4.189872e-27, 4.165455e-27, 4.169873e-27, 
    4.187818e-27, 4.229218e-27, 4.215059e-27, 4.250858e-27, 4.250049e-27, 
    4.290404e-27, 4.272043e-27, 4.340781e-27, 4.321177e-27, 4.378015e-27, 
    4.36367e-27, 4.377336e-27, 4.373193e-27, 4.37739e-27, 4.356365e-27, 
    4.365363e-27, 4.346902e-27, 4.275472e-27, 4.296375e-27, 4.23474e-27, 
    4.198303e-27, 4.174532e-27, 4.157812e-27, 4.160173e-27, 4.164671e-27, 
    4.187923e-27, 4.210064e-27, 4.227145e-27, 4.238611e-27, 4.249932e-27, 
    4.28445e-27, 4.303019e-27, 4.344739e-27, 4.337213e-27, 4.349986e-27, 
    4.362246e-27, 4.382848e-27, 4.379456e-27, 4.388543e-27, 4.349666e-27, 
    4.375469e-27, 4.332925e-27, 4.34453e-27, 4.25292e-27, 4.21888e-27, 
    4.204475e-27, 4.192026e-27, 4.161987e-27, 4.182645e-27, 4.174491e-27, 
    4.194043e-27, 4.206539e-27, 4.200359e-27, 4.238924e-27, 4.223847e-27, 
    4.304121e-27, 4.269147e-27, 4.360815e-27, 4.338759e-27, 4.366116e-27, 
    4.352147e-27, 4.376092e-27, 4.354538e-27, 4.391936e-27, 4.400098e-27, 
    4.394518e-27, 4.416011e-27, 4.353342e-27, 4.377327e-27, 4.200182e-27, 
    4.201189e-27, 4.205892e-27, 4.185241e-27, 4.183985e-27, 4.16533e-27, 
    4.181922e-27, 4.18906e-27, 4.207271e-27, 4.218115e-27, 4.228501e-27, 
    4.251398e-27, 4.277147e-27, 4.313748e-27, 4.340186e-27, 4.357964e-27, 
    4.347063e-27, 4.356686e-27, 4.345926e-27, 4.340894e-27, 4.397032e-27, 
    4.365442e-27, 4.412915e-27, 4.410283e-27, 4.388756e-27, 4.410579e-27, 
    4.201897e-27, 4.196102e-27, 4.17606e-27, 4.191725e-27, 4.163304e-27, 
    4.179132e-27, 4.188304e-27, 4.224142e-27, 4.232125e-27, 4.239507e-27, 
    4.254135e-27, 4.272981e-27, 4.306591e-27, 4.335992e-27, 4.362964e-27, 
    4.360985e-27, 4.361681e-27, 4.367711e-27, 4.352772e-27, 4.370167e-27, 
    4.373082e-27, 4.365449e-27, 4.40993e-27, 4.397192e-27, 4.410227e-27, 
    4.401932e-27, 4.197987e-27, 4.207749e-27, 4.202471e-27, 4.212396e-27, 
    4.205395e-27, 4.236829e-27, 4.246307e-27, 4.29117e-27, 4.272599e-27, 
    4.302209e-27, 4.275608e-27, 4.280307e-27, 4.303137e-27, 4.277048e-27, 
    4.334349e-27, 4.295412e-27, 4.367945e-27, 4.32882e-27, 4.370402e-27, 
    4.362846e-27, 4.375371e-27, 4.386598e-27, 4.400768e-27, 4.426966e-27, 
    4.420894e-27, 4.442878e-27, 4.222451e-27, 4.235299e-27, 4.234184e-27, 
    4.247668e-27, 4.257655e-27, 4.279504e-27, 4.314988e-27, 4.301628e-27, 
    4.326196e-27, 4.331133e-27, 4.293828e-27, 4.31669e-27, 4.243926e-27, 
    4.255502e-27, 4.24862e-27, 4.223454e-27, 4.30468e-27, 4.262616e-27, 
    4.34062e-27, 4.317613e-27, 4.384994e-27, 4.351378e-27, 4.41755e-27, 
    4.445995e-27, 4.472964e-27, 4.504519e-27, 4.242341e-27, 4.233597e-27, 
    4.249279e-27, 4.271015e-27, 4.291588e-27, 4.319011e-27, 4.321833e-27, 
    4.326981e-27, 4.340355e-27, 4.351613e-27, 4.328592e-27, 4.35444e-27, 
    4.258154e-27, 4.308362e-27, 4.230278e-27, 4.253504e-27, 4.269732e-27, 
    4.262626e-27, 4.300108e-27, 4.308994e-27, 4.345226e-27, 4.326481e-27, 
    4.438947e-27, 4.388947e-27, 4.528706e-27, 4.489342e-27, 4.23054e-27, 
    4.242319e-27, 4.28365e-27, 4.263856e-27, 4.320855e-27, 4.334979e-27, 
    4.346499e-27, 4.361226e-27, 4.362831e-27, 4.371577e-27, 4.357249e-27, 
    4.371017e-27, 4.319069e-27, 4.342235e-27, 4.278886e-27, 4.294239e-27, 
    4.287176e-27, 4.279428e-27, 4.303372e-27, 4.328949e-27, 4.329525e-27, 
    4.337744e-27, 4.360909e-27, 4.321088e-27, 4.445374e-27, 4.368289e-27, 
    4.255188e-27, 4.278054e-27, 4.281393e-27, 4.272429e-27, 4.33356e-27, 
    4.31134e-27, 4.371368e-27, 4.355095e-27, 4.381786e-27, 4.368507e-27, 
    4.366554e-27, 4.34955e-27, 4.338978e-27, 4.312352e-27, 4.290774e-27, 
    4.273732e-27, 4.277693e-27, 4.296431e-27, 4.330524e-27, 4.362964e-27, 
    4.35584e-27, 4.379755e-27, 4.316697e-27, 4.343048e-27, 4.332842e-27, 
    4.359495e-27, 4.301268e-27, 4.350731e-27, 4.288672e-27, 4.294098e-27, 
    4.3109e-27, 4.34482e-27, 4.352392e-27, 4.360434e-27, 4.355476e-27, 
    4.331397e-27, 4.327473e-27, 4.310498e-27, 4.305805e-27, 4.292919e-27, 
    4.282254e-27, 4.291991e-27, 4.302223e-27, 4.331419e-27, 4.357827e-27, 
    4.386754e-27, 4.393864e-27, 4.427788e-27, 4.400119e-27, 4.445801e-27, 
    4.406882e-27, 4.474428e-27, 4.353652e-27, 4.4058e-27, 4.311675e-27, 
    4.321757e-27, 4.340001e-27, 4.382103e-27, 4.35937e-27, 4.385978e-27, 
    4.327322e-27, 4.297064e-27, 4.289291e-27, 4.274761e-27, 4.289623e-27, 
    4.288415e-27, 4.302667e-27, 4.298087e-27, 4.332391e-27, 4.313942e-27, 
    4.366497e-27, 4.385775e-27, 4.44056e-27, 4.474353e-27, 4.508975e-27, 
    4.524301e-27, 4.528976e-27, 4.530929e-27,
  2.173993e-32, 2.192369e-32, 2.18878e-32, 2.203723e-32, 2.195421e-32, 
    2.205241e-32, 2.177705e-32, 2.193097e-32, 2.183247e-32, 2.175646e-32, 
    2.233275e-32, 2.2044e-32, 2.264059e-32, 2.245033e-32, 2.293091e-32, 
    2.261082e-32, 2.299593e-32, 2.292177e-32, 2.31459e-32, 2.308152e-32, 
    2.336984e-32, 2.317567e-32, 2.352068e-32, 2.332342e-32, 2.335414e-32, 
    2.316926e-32, 2.2102e-32, 2.229659e-32, 2.209048e-32, 2.211814e-32, 
    2.210576e-32, 2.195587e-32, 2.188108e-32, 2.172606e-32, 2.175412e-32, 
    2.186805e-32, 2.213059e-32, 2.204061e-32, 2.226823e-32, 2.226307e-32, 
    2.252035e-32, 2.240314e-32, 2.284413e-32, 2.271797e-32, 2.308421e-32, 
    2.299163e-32, 2.307983e-32, 2.305307e-32, 2.308018e-32, 2.294454e-32, 
    2.300256e-32, 2.288355e-32, 2.242488e-32, 2.255867e-32, 2.216569e-32, 
    2.193447e-32, 2.178374e-32, 2.167754e-32, 2.169253e-32, 2.172109e-32, 
    2.186872e-32, 2.200892e-32, 2.211739e-32, 2.219029e-32, 2.226232e-32, 
    2.248224e-32, 2.260134e-32, 2.286964e-32, 2.282115e-32, 2.290344e-32, 
    2.298245e-32, 2.311543e-32, 2.309352e-32, 2.315223e-32, 2.290135e-32, 
    2.306779e-32, 2.279354e-32, 2.286827e-32, 2.228148e-32, 2.206488e-32, 
    2.197356e-32, 2.189468e-32, 2.170405e-32, 2.183532e-32, 2.178348e-32, 
    2.190743e-32, 2.198658e-32, 2.194742e-32, 2.219229e-32, 2.209644e-32, 
    2.260842e-32, 2.238476e-32, 2.297322e-32, 2.283111e-32, 2.300741e-32, 
    2.291733e-32, 2.307181e-32, 2.293274e-32, 2.317415e-32, 2.322693e-32, 
    2.319084e-32, 2.33299e-32, 2.292504e-32, 2.307978e-32, 2.194631e-32, 
    2.195268e-32, 2.198248e-32, 2.185174e-32, 2.184379e-32, 2.172527e-32, 
    2.183071e-32, 2.18759e-32, 2.199121e-32, 2.206002e-32, 2.212601e-32, 
    2.227167e-32, 2.243551e-32, 2.267025e-32, 2.284029e-32, 2.295483e-32, 
    2.288457e-32, 2.294659e-32, 2.287725e-32, 2.284483e-32, 2.320711e-32, 
    2.300308e-32, 2.330985e-32, 2.329281e-32, 2.315361e-32, 2.329473e-32, 
    2.195717e-32, 2.192046e-32, 2.179345e-32, 2.189275e-32, 2.17124e-32, 
    2.181298e-32, 2.187114e-32, 2.209834e-32, 2.214905e-32, 2.2196e-32, 
    2.228909e-32, 2.240908e-32, 2.262426e-32, 2.281331e-32, 2.298707e-32, 
    2.297431e-32, 2.29788e-32, 2.30177e-32, 2.292137e-32, 2.303355e-32, 
    2.305238e-32, 2.300311e-32, 2.329052e-32, 2.320812e-32, 2.329244e-32, 
    2.323877e-32, 2.19324e-32, 2.199425e-32, 2.19608e-32, 2.202371e-32, 
    2.197934e-32, 2.217899e-32, 2.22393e-32, 2.25253e-32, 2.240667e-32, 
    2.259612e-32, 2.242573e-32, 2.24556e-32, 2.260214e-32, 2.243485e-32, 
    2.280276e-32, 2.255252e-32, 2.301921e-32, 2.276721e-32, 2.303507e-32, 
    2.298631e-32, 2.306713e-32, 2.313965e-32, 2.323125e-32, 2.340088e-32, 
    2.336153e-32, 2.350405e-32, 2.208756e-32, 2.216925e-32, 2.216214e-32, 
    2.224792e-32, 2.231152e-32, 2.245044e-32, 2.26782e-32, 2.259237e-32, 
    2.275025e-32, 2.278202e-32, 2.254229e-32, 2.268915e-32, 2.222412e-32, 
    2.229784e-32, 2.225399e-32, 2.209395e-32, 2.2612e-32, 2.234316e-32, 
    2.284309e-32, 2.269507e-32, 2.312929e-32, 2.291242e-32, 2.333987e-32, 
    2.352434e-32, 2.369946e-32, 2.390496e-32, 2.221403e-32, 2.21584e-32, 
    2.225817e-32, 2.239666e-32, 2.252793e-32, 2.270406e-32, 2.272219e-32, 
    2.27553e-32, 2.284137e-32, 2.29139e-32, 2.27657e-32, 2.293211e-32, 
    2.231479e-32, 2.263564e-32, 2.213732e-32, 2.228512e-32, 2.238849e-32, 
    2.234319e-32, 2.25826e-32, 2.263967e-32, 2.287277e-32, 2.275208e-32, 
    2.347862e-32, 2.315487e-32, 2.406272e-32, 2.380608e-32, 2.213897e-32, 
    2.221388e-32, 2.247704e-32, 2.235102e-32, 2.27159e-32, 2.280677e-32, 
    2.288094e-32, 2.297588e-32, 2.298622e-32, 2.304266e-32, 2.295022e-32, 
    2.303904e-32, 2.270443e-32, 2.285348e-32, 2.24465e-32, 2.254494e-32, 
    2.249962e-32, 2.244994e-32, 2.260356e-32, 2.2768e-32, 2.277167e-32, 
    2.282458e-32, 2.297398e-32, 2.27174e-32, 2.35204e-32, 2.302156e-32, 
    2.229579e-32, 2.244128e-32, 2.246256e-32, 2.240558e-32, 2.279764e-32, 
    2.265475e-32, 2.30413e-32, 2.293634e-32, 2.310856e-32, 2.302284e-32, 
    2.301024e-32, 2.29006e-32, 2.283252e-32, 2.266126e-32, 2.252273e-32, 
    2.241383e-32, 2.243893e-32, 2.255902e-32, 2.277812e-32, 2.298709e-32, 
    2.294116e-32, 2.309544e-32, 2.268917e-32, 2.285874e-32, 2.279303e-32, 
    2.296471e-32, 2.259006e-32, 2.290834e-32, 2.250922e-32, 2.254403e-32, 
    2.265193e-32, 2.287018e-32, 2.291891e-32, 2.297078e-32, 2.293879e-32, 
    2.278374e-32, 2.275848e-32, 2.264933e-32, 2.26192e-32, 2.253646e-32, 
    2.246806e-32, 2.253051e-32, 2.259621e-32, 2.278386e-32, 2.295397e-32, 
    2.314067e-32, 2.31866e-32, 2.340628e-32, 2.322712e-32, 2.352317e-32, 
    2.327098e-32, 2.37091e-32, 2.292711e-32, 2.326389e-32, 2.265689e-32, 
    2.27217e-32, 2.283914e-32, 2.311066e-32, 2.29639e-32, 2.313568e-32, 
    2.27575e-32, 2.25631e-32, 2.25132e-32, 2.242036e-32, 2.251533e-32, 
    2.250757e-32, 2.259903e-32, 2.256962e-32, 2.279011e-32, 2.267146e-32, 
    2.300988e-32, 2.313436e-32, 2.348903e-32, 2.370854e-32, 2.393396e-32, 
    2.403395e-32, 2.406446e-32, 2.407722e-32,
  3.734964e-38, 3.774637e-38, 3.766887e-38, 3.79918e-38, 3.78123e-38, 
    3.80245e-38, 3.742974e-38, 3.776215e-38, 3.754949e-38, 3.738528e-38, 
    3.863047e-38, 3.800639e-38, 3.92982e-38, 3.888498e-38, 3.993215e-38, 
    3.923346e-38, 4.007596e-38, 3.991204e-38, 4.040998e-38, 4.02664e-38, 
    4.091139e-38, 4.047643e-38, 4.125064e-38, 4.080717e-38, 4.087611e-38, 
    4.046213e-38, 3.813135e-38, 3.855212e-38, 3.810652e-38, 3.81662e-38, 
    3.813946e-38, 3.781592e-38, 3.765443e-38, 3.731967e-38, 3.738022e-38, 
    3.762627e-38, 3.819307e-38, 3.799903e-38, 3.849046e-38, 3.84793e-38, 
    3.903682e-38, 3.878287e-38, 3.974213e-38, 3.946666e-38, 4.027238e-38, 
    4.006634e-38, 4.026264e-38, 4.020303e-38, 4.026341e-38, 3.996193e-38, 
    4.009066e-38, 3.982834e-38, 3.88299e-38, 3.912003e-38, 3.826882e-38, 
    3.776977e-38, 3.744419e-38, 3.721507e-38, 3.724738e-38, 3.7309e-38, 
    3.762772e-38, 3.793064e-38, 3.816452e-38, 3.832192e-38, 3.847769e-38, 
    3.895428e-38, 3.921283e-38, 3.979797e-38, 3.969188e-38, 3.987193e-38, 
    4.004592e-38, 4.034201e-38, 4.029314e-38, 4.042413e-38, 3.986731e-38, 
    4.023586e-38, 3.963154e-38, 3.979491e-38, 3.85194e-38, 3.805131e-38, 
    3.785425e-38, 3.768373e-38, 3.727222e-38, 3.755567e-38, 3.744365e-38, 
    3.771121e-38, 3.78823e-38, 3.779762e-38, 3.832623e-38, 3.811934e-38, 
    3.922821e-38, 3.874311e-38, 4.002542e-38, 3.971364e-38, 4.010141e-38, 
    3.990229e-38, 4.024479e-38, 3.993606e-38, 4.047306e-38, 4.059108e-38, 
    4.051037e-38, 4.082163e-38, 3.991919e-38, 4.026256e-38, 3.779521e-38, 
    3.7809e-38, 3.787342e-38, 3.75911e-38, 3.757394e-38, 3.731798e-38, 
    3.754567e-38, 3.76432e-38, 3.78923e-38, 3.804085e-38, 3.818314e-38, 
    3.849795e-38, 3.885293e-38, 3.936273e-38, 3.973373e-38, 3.998454e-38, 
    3.983057e-38, 3.99664e-38, 3.981456e-38, 3.974364e-38, 4.054676e-38, 
    4.009182e-38, 4.07767e-38, 4.073849e-38, 4.042722e-38, 4.07428e-38, 
    3.78187e-38, 3.773936e-38, 3.746516e-38, 3.767953e-38, 3.729023e-38, 
    3.750738e-38, 3.763295e-38, 3.812349e-38, 3.823284e-38, 3.833429e-38, 
    3.853565e-38, 3.879572e-38, 3.926263e-38, 3.967478e-38, 4.005618e-38, 
    4.002782e-38, 4.003779e-38, 4.012431e-38, 3.991115e-38, 4.015958e-38, 
    4.020152e-38, 4.009186e-38, 4.073337e-38, 4.054896e-38, 4.073768e-38, 
    4.061751e-38, 3.776515e-38, 3.789889e-38, 3.782655e-38, 3.796266e-38, 
    3.786666e-38, 3.829759e-38, 3.842798e-38, 3.904762e-38, 3.879053e-38, 
    3.920144e-38, 3.883172e-38, 3.88964e-38, 3.921464e-38, 3.885144e-38, 
    3.965179e-38, 3.910676e-38, 4.012768e-38, 3.957422e-38, 4.016296e-38, 
    4.00545e-38, 4.023433e-38, 4.039606e-38, 4.060068e-38, 4.098103e-38, 
    4.089264e-38, 4.121312e-38, 3.81002e-38, 3.827652e-38, 3.82611e-38, 
    3.844654e-38, 3.858425e-38, 3.888518e-38, 3.938003e-38, 3.919322e-38, 
    3.953705e-38, 3.960641e-38, 3.908441e-38, 3.94039e-38, 3.839509e-38, 
    3.855468e-38, 3.845968e-38, 3.8114e-38, 3.923598e-38, 3.865288e-38, 
    3.973986e-38, 3.941676e-38, 4.037294e-38, 3.989161e-38, 4.084403e-38, 
    4.125896e-38, 4.16545e-38, 4.212139e-38, 3.837325e-38, 3.825303e-38, 
    3.846869e-38, 3.876893e-38, 3.905327e-38, 3.943636e-38, 3.947586e-38, 
    3.95481e-38, 3.973607e-38, 3.989477e-38, 3.957083e-38, 3.993468e-38, 
    3.85915e-38, 3.928739e-38, 3.820755e-38, 3.852715e-38, 3.87512e-38, 
    3.865289e-38, 3.917196e-38, 3.92961e-38, 3.98048e-38, 3.954104e-38, 
    4.115599e-38, 4.04301e-38, 4.248142e-38, 4.189643e-38, 3.821108e-38, 
    3.83729e-38, 3.89429e-38, 3.866988e-38, 3.946215e-38, 3.966048e-38, 
    3.982262e-38, 4.003136e-38, 4.00543e-38, 4.017987e-38, 3.997436e-38, 
    4.017178e-38, 3.943718e-38, 3.976257e-38, 3.887663e-38, 3.90902e-38, 
    3.899181e-38, 3.888409e-38, 3.921754e-38, 3.957587e-38, 3.95838e-38, 
    3.969942e-38, 4.002741e-38, 3.946541e-38, 4.125029e-38, 4.013317e-38, 
    3.855016e-38, 3.886543e-38, 3.891145e-38, 3.878813e-38, 3.964054e-38, 
    3.932895e-38, 4.017684e-38, 3.994393e-38, 4.032667e-38, 4.013573e-38, 
    4.010772e-38, 3.986566e-38, 3.971673e-38, 3.934314e-38, 3.904198e-38, 
    3.880596e-38, 3.886026e-38, 3.912078e-38, 3.959796e-38, 4.005627e-38, 
    3.995457e-38, 4.029741e-38, 3.94039e-38, 3.97741e-38, 3.96305e-38, 
    4.00065e-38, 3.918821e-38, 3.988287e-38, 3.901263e-38, 3.908818e-38, 
    3.93228e-38, 3.979919e-38, 3.990576e-38, 4.002001e-38, 3.994932e-38, 
    3.96102e-38, 3.955504e-38, 3.931714e-38, 3.92516e-38, 3.907174e-38, 
    3.892336e-38, 3.905885e-38, 3.92016e-38, 3.961044e-38, 3.998268e-38, 
    4.039833e-38, 4.050086e-38, 4.099332e-38, 4.059161e-38, 4.125656e-38, 
    4.068997e-38, 4.167661e-38, 3.992387e-38, 4.067392e-38, 3.933359e-38, 
    3.947478e-38, 3.973127e-38, 4.033148e-38, 4.000471e-38, 4.038727e-38, 
    3.95529e-38, 3.91297e-38, 3.902126e-38, 3.88201e-38, 3.902589e-38, 
    3.900906e-38, 3.920769e-38, 3.914376e-38, 3.962409e-38, 3.936532e-38, 
    4.010695e-38, 4.038429e-38, 4.117932e-38, 4.167518e-38, 4.218731e-38, 
    4.241557e-38, 4.248535e-38, 4.251455e-38,
  2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.522337e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.662467e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  2.094773e-05, 2.075879e-05, 2.079557e-05, 2.064283e-05, 2.072761e-05, 
    2.062752e-05, 2.090948e-05, 2.075127e-05, 2.085232e-05, 2.093075e-05, 
    2.034529e-05, 2.063601e-05, 2.004194e-05, 2.02284e-05, 1.975899e-05, 
    2.007098e-05, 1.969591e-05, 1.976804e-05, 1.955076e-05, 1.961308e-05, 
    1.933434e-05, 1.952197e-05, 1.918943e-05, 1.937921e-05, 1.934955e-05, 
    1.952815e-05, 2.057763e-05, 2.038155e-05, 2.058922e-05, 2.056131e-05, 
    2.057384e-05, 2.072585e-05, 2.08023e-05, 2.096215e-05, 2.093317e-05, 
    2.081575e-05, 2.054875e-05, 2.063953e-05, 2.041052e-05, 2.04157e-05, 
    2.015975e-05, 2.027529e-05, 1.984355e-05, 1.996656e-05, 1.961048e-05, 
    1.970021e-05, 1.961469e-05, 1.964064e-05, 1.961435e-05, 1.97459e-05, 
    1.968957e-05, 1.980522e-05, 2.025366e-05, 2.012219e-05, 2.051347e-05, 
    2.074753e-05, 2.090254e-05, 2.101228e-05, 2.099678e-05, 2.096721e-05, 
    2.081507e-05, 2.067168e-05, 2.056218e-05, 2.048881e-05, 2.041645e-05, 
    2.019683e-05, 2.008032e-05, 1.981864e-05, 1.986596e-05, 1.978579e-05, 
    1.970913e-05, 1.95802e-05, 1.960144e-05, 1.954457e-05, 1.978792e-05, 
    1.962628e-05, 1.989289e-05, 1.982008e-05, 2.039669e-05, 2.061506e-05, 
    2.070758e-05, 2.07885e-05, 2.098486e-05, 2.084932e-05, 2.090279e-05, 
    2.077552e-05, 2.069451e-05, 2.073459e-05, 2.048681e-05, 2.058326e-05, 
    2.007341e-05, 2.029353e-05, 1.971807e-05, 1.985625e-05, 1.968491e-05, 
    1.97724e-05, 1.962242e-05, 1.975742e-05, 1.95234e-05, 1.947233e-05, 
    1.950723e-05, 1.937307e-05, 1.976489e-05, 1.961469e-05, 2.073571e-05, 
    2.072918e-05, 2.069873e-05, 2.083247e-05, 2.084064e-05, 2.096295e-05, 
    2.085414e-05, 2.080774e-05, 2.068982e-05, 2.061994e-05, 2.055345e-05, 
    2.040701e-05, 2.024303e-05, 2.001304e-05, 1.98473e-05, 1.973596e-05, 
    1.980426e-05, 1.974397e-05, 1.981136e-05, 1.984293e-05, 1.949147e-05, 
    1.968904e-05, 1.939239e-05, 1.940884e-05, 1.954322e-05, 1.940699e-05, 
    2.072459e-05, 2.076219e-05, 2.089254e-05, 2.079056e-05, 2.097625e-05, 
    2.087237e-05, 2.081255e-05, 2.058123e-05, 2.05303e-05, 2.048302e-05, 
    2.038955e-05, 2.026938e-05, 2.0058e-05, 1.987353e-05, 1.970467e-05, 
    1.971706e-05, 1.97127e-05, 1.967491e-05, 1.976845e-05, 1.965954e-05, 
    1.964124e-05, 1.968908e-05, 1.941104e-05, 1.949059e-05, 1.940919e-05, 
    1.9461e-05, 2.074997e-05, 2.068668e-05, 2.072089e-05, 2.065654e-05, 
    2.070187e-05, 2.050001e-05, 2.043936e-05, 2.015477e-05, 2.027174e-05, 
    2.00855e-05, 2.025285e-05, 2.022323e-05, 2.007939e-05, 2.024382e-05, 
    1.98837e-05, 2.012805e-05, 1.967344e-05, 1.991823e-05, 1.965807e-05, 
    1.97054e-05, 1.962703e-05, 1.955675e-05, 1.946825e-05, 1.930461e-05, 
    1.934254e-05, 1.920548e-05, 2.05922e-05, 2.050987e-05, 2.051714e-05, 
    2.043088e-05, 2.036701e-05, 2.022836e-05, 2.000533e-05, 2.00893e-05, 
    1.993508e-05, 1.990407e-05, 2.013834e-05, 1.999459e-05, 2.045472e-05, 
    2.03806e-05, 2.042475e-05, 2.05857e-05, 2.006994e-05, 2.033516e-05, 
    1.984456e-05, 1.998888e-05, 1.956677e-05, 1.977703e-05, 1.936341e-05, 
    1.918577e-05, 1.901824e-05, 1.882186e-05, 2.046491e-05, 2.05209e-05, 
    2.042062e-05, 2.028159e-05, 2.015234e-05, 1.998009e-05, 1.996244e-05, 
    1.993011e-05, 1.984629e-05, 1.977573e-05, 1.991987e-05, 1.975803e-05, 
    2.036337e-05, 2.004687e-05, 2.054205e-05, 2.039334e-05, 2.02898e-05, 
    2.033525e-05, 2.009889e-05, 2.004305e-05, 1.981562e-05, 1.99333e-05, 
    1.922965e-05, 1.954188e-05, 1.867202e-05, 1.89162e-05, 2.054045e-05, 
    2.046511e-05, 2.020216e-05, 2.032741e-05, 1.996858e-05, 1.987994e-05, 
    1.98078e-05, 1.971544e-05, 1.970548e-05, 1.965069e-05, 1.974044e-05, 
    1.965424e-05, 1.997972e-05, 1.983447e-05, 2.023228e-05, 2.013568e-05, 
    2.018014e-05, 2.022887e-05, 2.007836e-05, 1.99176e-05, 1.991418e-05, 
    1.986254e-05, 1.971676e-05, 1.996712e-05, 1.91892e-05, 1.967067e-05, 
    2.038285e-05, 2.023724e-05, 2.021644e-05, 2.02729e-05, 1.988883e-05, 
    2.002826e-05, 1.965203e-05, 1.975393e-05, 1.958689e-05, 1.966995e-05, 
    1.968215e-05, 1.978866e-05, 1.985488e-05, 2.002187e-05, 2.015742e-05, 
    2.026472e-05, 2.023979e-05, 2.012187e-05, 1.990776e-05, 1.970456e-05, 
    1.974913e-05, 1.95996e-05, 1.999466e-05, 1.982929e-05, 1.989325e-05, 
    1.972634e-05, 2.009152e-05, 1.978062e-05, 2.017074e-05, 2.013663e-05, 
    2.003102e-05, 1.981804e-05, 1.977086e-05, 1.97204e-05, 1.975154e-05, 
    1.990232e-05, 1.992699e-05, 2.00336e-05, 2.006299e-05, 2.014406e-05, 
    2.02111e-05, 2.014985e-05, 2.008546e-05, 1.990226e-05, 1.973671e-05, 
    1.955575e-05, 1.951139e-05, 1.929914e-05, 1.947195e-05, 1.918651e-05, 
    1.942922e-05, 1.900856e-05, 1.976259e-05, 1.943638e-05, 2.002622e-05, 
    1.996294e-05, 1.984829e-05, 1.958464e-05, 1.972713e-05, 1.956046e-05, 
    1.992796e-05, 2.011779e-05, 2.016683e-05, 2.02582e-05, 2.016474e-05, 
    2.017235e-05, 2.00828e-05, 2.011159e-05, 1.989617e-05, 2.001198e-05, 
    1.968246e-05, 1.956178e-05, 1.921985e-05, 1.900937e-05, 1.879449e-05, 
    1.869941e-05, 1.867045e-05, 1.865833e-05,
  1.394598e-05, 1.376952e-05, 1.380386e-05, 1.366133e-05, 1.374043e-05, 
    1.364705e-05, 1.391024e-05, 1.37625e-05, 1.385685e-05, 1.393012e-05, 
    1.338408e-05, 1.365497e-05, 1.310205e-05, 1.327535e-05, 1.283952e-05, 
    1.312902e-05, 1.278106e-05, 1.284791e-05, 1.264668e-05, 1.270436e-05, 
    1.244658e-05, 1.262005e-05, 1.23128e-05, 1.248804e-05, 1.246063e-05, 
    1.262576e-05, 1.360054e-05, 1.341784e-05, 1.361135e-05, 1.358532e-05, 
    1.359701e-05, 1.373879e-05, 1.381014e-05, 1.395947e-05, 1.393238e-05, 
    1.38227e-05, 1.357361e-05, 1.365826e-05, 1.344484e-05, 1.344967e-05, 
    1.321152e-05, 1.331897e-05, 1.291792e-05, 1.303206e-05, 1.270196e-05, 
    1.278506e-05, 1.270586e-05, 1.272988e-05, 1.270554e-05, 1.28274e-05, 
    1.27752e-05, 1.288238e-05, 1.329885e-05, 1.317661e-05, 1.354074e-05, 
    1.375901e-05, 1.390376e-05, 1.400632e-05, 1.399183e-05, 1.396419e-05, 
    1.382206e-05, 1.368825e-05, 1.358614e-05, 1.351777e-05, 1.345036e-05, 
    1.324597e-05, 1.31377e-05, 1.289482e-05, 1.293871e-05, 1.286436e-05, 
    1.279332e-05, 1.267393e-05, 1.269359e-05, 1.264096e-05, 1.286634e-05, 
    1.271659e-05, 1.29637e-05, 1.289616e-05, 1.343193e-05, 1.363544e-05, 
    1.372172e-05, 1.379726e-05, 1.398068e-05, 1.385405e-05, 1.390399e-05, 
    1.378515e-05, 1.370955e-05, 1.374695e-05, 1.35159e-05, 1.360579e-05, 
    1.313127e-05, 1.333594e-05, 1.280161e-05, 1.292971e-05, 1.277089e-05, 
    1.285196e-05, 1.271301e-05, 1.283807e-05, 1.262137e-05, 1.257412e-05, 
    1.260641e-05, 1.248238e-05, 1.2845e-05, 1.270585e-05, 1.374799e-05, 
    1.374189e-05, 1.371348e-05, 1.383831e-05, 1.384594e-05, 1.396021e-05, 
    1.385855e-05, 1.381522e-05, 1.370517e-05, 1.363999e-05, 1.3578e-05, 
    1.344157e-05, 1.328896e-05, 1.307521e-05, 1.29214e-05, 1.281819e-05, 
    1.28815e-05, 1.28256e-05, 1.288808e-05, 1.291735e-05, 1.259182e-05, 
    1.277471e-05, 1.250022e-05, 1.251543e-05, 1.26397e-05, 1.251372e-05, 
    1.373761e-05, 1.377271e-05, 1.389442e-05, 1.379918e-05, 1.397264e-05, 
    1.387558e-05, 1.381971e-05, 1.360389e-05, 1.355643e-05, 1.351237e-05, 
    1.342531e-05, 1.331347e-05, 1.311697e-05, 1.294572e-05, 1.278919e-05, 
    1.280067e-05, 1.279663e-05, 1.276162e-05, 1.28483e-05, 1.274739e-05, 
    1.273044e-05, 1.277474e-05, 1.251746e-05, 1.259102e-05, 1.251575e-05, 
    1.256365e-05, 1.37613e-05, 1.370224e-05, 1.373416e-05, 1.367412e-05, 
    1.371642e-05, 1.352819e-05, 1.347168e-05, 1.320689e-05, 1.331567e-05, 
    1.314251e-05, 1.32981e-05, 1.327054e-05, 1.313682e-05, 1.32897e-05, 
    1.295516e-05, 1.318204e-05, 1.276026e-05, 1.298718e-05, 1.274603e-05, 
    1.278987e-05, 1.271728e-05, 1.265223e-05, 1.257035e-05, 1.241912e-05, 
    1.245416e-05, 1.232761e-05, 1.361413e-05, 1.353739e-05, 1.354416e-05, 
    1.34638e-05, 1.340433e-05, 1.327532e-05, 1.306805e-05, 1.314605e-05, 
    1.300284e-05, 1.297406e-05, 1.319162e-05, 1.305808e-05, 1.3486e-05, 
    1.341697e-05, 1.345809e-05, 1.360807e-05, 1.312805e-05, 1.337467e-05, 
    1.291886e-05, 1.305279e-05, 1.26615e-05, 1.285624e-05, 1.247344e-05, 
    1.230942e-05, 1.215497e-05, 1.197418e-05, 1.34955e-05, 1.354767e-05, 
    1.345425e-05, 1.332482e-05, 1.320463e-05, 1.304462e-05, 1.302824e-05, 
    1.299823e-05, 1.292047e-05, 1.285505e-05, 1.298872e-05, 1.283864e-05, 
    1.340092e-05, 1.310663e-05, 1.356737e-05, 1.342883e-05, 1.333246e-05, 
    1.337476e-05, 1.315496e-05, 1.310308e-05, 1.289202e-05, 1.300119e-05, 
    1.23499e-05, 1.263845e-05, 1.183647e-05, 1.206098e-05, 1.356589e-05, 
    1.349568e-05, 1.325094e-05, 1.336747e-05, 1.303394e-05, 1.295167e-05, 
    1.288477e-05, 1.279917e-05, 1.278994e-05, 1.273919e-05, 1.282234e-05, 
    1.274248e-05, 1.304428e-05, 1.290951e-05, 1.327897e-05, 1.318915e-05, 
    1.323049e-05, 1.32758e-05, 1.313589e-05, 1.298661e-05, 1.298345e-05, 
    1.293553e-05, 1.280036e-05, 1.303258e-05, 1.231256e-05, 1.275766e-05, 
    1.341907e-05, 1.328357e-05, 1.326424e-05, 1.331675e-05, 1.295992e-05, 
    1.308935e-05, 1.274043e-05, 1.283484e-05, 1.268012e-05, 1.275702e-05, 
    1.276833e-05, 1.286703e-05, 1.292843e-05, 1.308341e-05, 1.320936e-05, 
    1.330914e-05, 1.328595e-05, 1.317631e-05, 1.297748e-05, 1.278909e-05, 
    1.283038e-05, 1.269189e-05, 1.305815e-05, 1.290469e-05, 1.296402e-05, 
    1.280927e-05, 1.314811e-05, 1.285954e-05, 1.322174e-05, 1.319004e-05, 
    1.309191e-05, 1.289426e-05, 1.285053e-05, 1.280376e-05, 1.283263e-05, 
    1.297243e-05, 1.299534e-05, 1.309431e-05, 1.31216e-05, 1.319694e-05, 
    1.325927e-05, 1.320232e-05, 1.314248e-05, 1.297239e-05, 1.281887e-05, 
    1.265129e-05, 1.261026e-05, 1.241405e-05, 1.257376e-05, 1.231007e-05, 
    1.253422e-05, 1.214602e-05, 1.284284e-05, 1.254087e-05, 1.308746e-05, 
    1.30287e-05, 1.292232e-05, 1.267802e-05, 1.281e-05, 1.265565e-05, 
    1.299624e-05, 1.317251e-05, 1.321811e-05, 1.330307e-05, 1.321617e-05, 
    1.322324e-05, 1.314002e-05, 1.316677e-05, 1.296674e-05, 1.307423e-05, 
    1.276861e-05, 1.265688e-05, 1.234087e-05, 1.214678e-05, 1.194903e-05, 
    1.186163e-05, 1.183503e-05, 1.18239e-05,
  5.604251e-06, 5.50667e-06, 5.525618e-06, 5.44709e-06, 5.49063e-06, 
    5.439244e-06, 5.584448e-06, 5.502797e-06, 5.554899e-06, 5.595462e-06, 
    5.295302e-06, 5.443593e-06, 5.142209e-06, 5.236123e-06, 5.000915e-06, 
    5.156791e-06, 4.969615e-06, 5.005412e-06, 4.897878e-06, 4.928632e-06, 
    4.791638e-06, 4.883699e-06, 4.721001e-06, 4.813595e-06, 4.799076e-06, 
    4.88674e-06, 5.4137e-06, 5.313715e-06, 5.419632e-06, 5.40535e-06, 
    5.411761e-06, 5.489725e-06, 5.529085e-06, 5.611732e-06, 5.596713e-06, 
    5.536025e-06, 5.39893e-06, 5.445404e-06, 5.328458e-06, 5.331093e-06, 
    5.201477e-06, 5.259838e-06, 5.04299e-06, 5.104429e-06, 4.927348e-06, 
    4.97175e-06, 4.929429e-06, 4.942255e-06, 4.929262e-06, 4.994419e-06, 
    4.966479e-06, 5.023903e-06, 5.248894e-06, 5.182551e-06, 5.380914e-06, 
    5.50087e-06, 5.58086e-06, 5.637738e-06, 5.629691e-06, 5.614353e-06, 
    5.53567e-06, 5.461896e-06, 5.405798e-06, 5.368334e-06, 5.331472e-06, 
    5.220169e-06, 5.161487e-06, 5.030579e-06, 5.054163e-06, 5.014234e-06, 
    4.976172e-06, 4.912398e-06, 4.922884e-06, 4.89483e-06, 5.015296e-06, 
    4.935156e-06, 5.067604e-06, 5.0313e-06, 5.321409e-06, 5.432861e-06, 
    5.480324e-06, 5.521973e-06, 5.623504e-06, 5.553349e-06, 5.580984e-06, 
    5.515292e-06, 5.473619e-06, 5.494224e-06, 5.36731e-06, 5.416581e-06, 
    5.158013e-06, 5.269073e-06, 4.980609e-06, 5.049321e-06, 4.964172e-06, 
    5.007585e-06, 4.933247e-06, 5.000139e-06, 4.884401e-06, 4.859275e-06, 
    4.876441e-06, 4.810593e-06, 5.003852e-06, 4.929424e-06, 5.494799e-06, 
    5.491437e-06, 5.475786e-06, 5.544649e-06, 5.548869e-06, 5.612141e-06, 
    5.55584e-06, 5.531893e-06, 5.471209e-06, 5.435365e-06, 5.401338e-06, 
    5.32667e-06, 5.243518e-06, 5.127712e-06, 5.04486e-06, 4.989486e-06, 
    5.023428e-06, 4.993459e-06, 5.026962e-06, 5.042684e-06, 4.868683e-06, 
    4.966215e-06, 4.820051e-06, 4.828114e-06, 4.894161e-06, 4.827206e-06, 
    5.489077e-06, 5.508427e-06, 5.575688e-06, 5.523037e-06, 5.61904e-06, 
    5.565258e-06, 5.534373e-06, 5.415539e-06, 5.389509e-06, 5.365378e-06, 
    5.317795e-06, 5.256847e-06, 5.150276e-06, 5.057935e-06, 4.973962e-06, 
    4.980106e-06, 4.977942e-06, 4.959217e-06, 5.005621e-06, 4.951608e-06, 
    4.942552e-06, 4.966233e-06, 4.829194e-06, 4.868257e-06, 4.828286e-06, 
    4.853712e-06, 5.502137e-06, 5.469597e-06, 5.487175e-06, 5.454126e-06, 
    5.477401e-06, 5.37404e-06, 5.343125e-06, 5.198962e-06, 5.258043e-06, 
    5.164095e-06, 5.248487e-06, 5.23351e-06, 5.161015e-06, 5.243923e-06, 
    5.063007e-06, 5.185498e-06, 4.95849e-06, 5.080245e-06, 4.95088e-06, 
    4.974325e-06, 4.935527e-06, 4.900832e-06, 4.857271e-06, 4.777116e-06, 
    4.795651e-06, 4.728806e-06, 5.421159e-06, 5.379076e-06, 5.382788e-06, 
    5.338818e-06, 5.306343e-06, 5.236106e-06, 5.123849e-06, 5.166005e-06, 
    5.088679e-06, 5.073182e-06, 5.190687e-06, 5.118464e-06, 5.350955e-06, 
    5.313241e-06, 5.335696e-06, 5.417831e-06, 5.156272e-06, 5.290172e-06, 
    5.043492e-06, 5.115608e-06, 4.905774e-06, 5.009877e-06, 4.80586e-06, 
    4.719219e-06, 4.638063e-06, 4.543608e-06, 5.356146e-06, 5.384708e-06, 
    5.333596e-06, 5.263023e-06, 5.197741e-06, 5.111201e-06, 5.102369e-06, 
    5.086194e-06, 5.04436e-06, 5.009239e-06, 5.081073e-06, 5.000445e-06, 
    5.304482e-06, 5.144687e-06, 5.395506e-06, 5.319713e-06, 5.267182e-06, 
    5.290222e-06, 5.170831e-06, 5.142771e-06, 5.029079e-06, 5.087788e-06, 
    4.74056e-06, 4.893497e-06, 4.472044e-06, 4.588888e-06, 5.394693e-06, 
    5.356249e-06, 5.222867e-06, 5.286247e-06, 5.10544e-06, 5.061135e-06, 
    5.025187e-06, 4.979303e-06, 4.974362e-06, 4.947226e-06, 4.991708e-06, 
    4.948985e-06, 5.111017e-06, 5.038469e-06, 5.23809e-06, 5.189348e-06, 
    5.211763e-06, 5.236365e-06, 5.16051e-06, 5.079938e-06, 5.078235e-06, 
    5.052456e-06, 4.97994e-06, 5.10471e-06, 4.720876e-06, 4.957101e-06, 
    5.314389e-06, 5.24059e-06, 5.230085e-06, 5.258632e-06, 5.065572e-06, 
    5.135347e-06, 4.947889e-06, 4.998406e-06, 4.9157e-06, 4.956758e-06, 
    4.962804e-06, 5.015666e-06, 5.048636e-06, 5.13214e-06, 5.200302e-06, 
    5.254492e-06, 5.241882e-06, 5.182392e-06, 5.075022e-06, 4.973907e-06, 
    4.996016e-06, 4.921975e-06, 5.118505e-06, 5.035883e-06, 5.067777e-06, 
    4.98471e-06, 5.167123e-06, 5.011652e-06, 5.207019e-06, 5.18983e-06, 
    5.136734e-06, 5.03028e-06, 5.006816e-06, 4.981761e-06, 4.997221e-06, 
    5.072305e-06, 5.084636e-06, 5.138027e-06, 5.152782e-06, 5.193572e-06, 
    5.227386e-06, 5.196486e-06, 5.164073e-06, 5.07228e-06, 4.989854e-06, 
    4.900336e-06, 4.87849e-06, 4.774435e-06, 4.85908e-06, 4.719564e-06, 
    4.838088e-06, 4.633377e-06, 5.002697e-06, 4.841614e-06, 5.134326e-06, 
    5.102616e-06, 5.04535e-06, 4.91458e-06, 4.985101e-06, 4.902657e-06, 
    5.085121e-06, 5.180334e-06, 5.205048e-06, 5.251191e-06, 5.203994e-06, 
    5.20783e-06, 5.162743e-06, 5.177224e-06, 5.069238e-06, 5.127184e-06, 
    4.962952e-06, 4.903311e-06, 4.735796e-06, 4.633777e-06, 4.53051e-06, 
    4.485096e-06, 4.471297e-06, 4.465531e-06,
  1.104519e-06, 1.075676e-06, 1.081255e-06, 1.058202e-06, 1.070961e-06, 
    1.055909e-06, 1.098643e-06, 1.074537e-06, 1.089896e-06, 1.101909e-06, 
    1.01416e-06, 1.05718e-06, 9.704301e-07, 9.971722e-07, 9.30695e-07, 
    9.745653e-07, 9.21974e-07, 9.3195e-07, 9.020992e-07, 9.106004e-07, 
    8.729549e-07, 8.981894e-07, 8.537688e-07, 8.789496e-07, 8.74984e-07, 
    8.990276e-07, 1.048455e-06, 1.019466e-06, 1.050185e-06, 1.046023e-06, 
    1.04789e-06, 1.070696e-06, 1.082277e-06, 1.106741e-06, 1.102281e-06, 
    1.084323e-06, 1.044154e-06, 1.057709e-06, 1.023721e-06, 1.024483e-06, 
    9.872758e-07, 1.003967e-06, 9.424641e-07, 9.59746e-07, 9.102449e-07, 
    9.225677e-07, 9.108211e-07, 9.143754e-07, 9.107749e-07, 9.288823e-07, 
    9.211017e-07, 9.371182e-07, 1.000829e-06, 9.818851e-07, 1.038917e-06, 
    1.073971e-06, 1.097579e-06, 1.11448e-06, 1.112084e-06, 1.10752e-06, 
    1.084219e-06, 1.062535e-06, 1.046153e-06, 1.035265e-06, 1.024592e-06, 
    9.926114e-07, 9.758979e-07, 9.389871e-07, 9.455983e-07, 9.344147e-07, 
    9.237984e-07, 9.061094e-07, 9.090094e-07, 9.012581e-07, 9.347113e-07, 
    9.124077e-07, 9.493738e-07, 9.391887e-07, 1.021687e-06, 1.054044e-06, 
    1.067937e-06, 1.080181e-06, 1.110242e-06, 1.089438e-06, 1.097616e-06, 
    1.078213e-06, 1.06597e-06, 1.072017e-06, 1.034968e-06, 1.049295e-06, 
    9.749118e-07, 1.006617e-06, 9.250335e-07, 9.442397e-07, 9.204603e-07, 
    9.325565e-07, 9.118787e-07, 9.304779e-07, 8.983831e-07, 8.914695e-07, 
    8.961908e-07, 8.781288e-07, 9.315143e-07, 9.1082e-07, 1.072186e-06, 
    1.071198e-06, 1.066605e-06, 1.086869e-06, 1.088115e-06, 1.106863e-06, 
    1.090175e-06, 1.083105e-06, 1.065263e-06, 1.054776e-06, 1.044855e-06, 
    1.023205e-06, 9.992893e-07, 9.663253e-07, 9.429884e-07, 9.275067e-07, 
    9.369853e-07, 9.286143e-07, 9.379741e-07, 9.42378e-07, 8.940559e-07, 
    9.210286e-07, 8.80715e-07, 8.82922e-07, 9.010737e-07, 8.826732e-07, 
    1.070505e-06, 1.076192e-06, 1.096047e-06, 1.080494e-06, 1.108914e-06, 
    1.09296e-06, 1.083836e-06, 1.048992e-06, 1.041414e-06, 1.034408e-06, 
    1.020642e-06, 1.003109e-06, 9.727166e-07, 9.466575e-07, 9.231833e-07, 
    9.248932e-07, 9.24291e-07, 9.190834e-07, 9.320083e-07, 9.169705e-07, 
    9.144576e-07, 9.210333e-07, 8.832177e-07, 8.939385e-07, 8.829689e-07, 
    8.89941e-07, 1.074342e-06, 1.064791e-06, 1.069947e-06, 1.06026e-06, 
    1.067079e-06, 1.036921e-06, 1.027962e-06, 9.865591e-07, 1.003452e-06, 
    9.766383e-07, 1.000712e-06, 9.964245e-07, 9.757642e-07, 9.994048e-07, 
    9.480825e-07, 9.827241e-07, 9.188814e-07, 9.529305e-07, 9.167684e-07, 
    9.232841e-07, 9.125102e-07, 9.029145e-07, 8.909187e-07, 8.689977e-07, 
    8.740492e-07, 8.55881e-07, 1.05063e-06, 1.038383e-06, 1.039461e-06, 
    1.026716e-06, 1.01734e-06, 9.971671e-07, 9.652324e-07, 9.771808e-07, 
    9.553049e-07, 9.509425e-07, 9.842009e-07, 9.637102e-07, 1.030228e-06, 
    1.019329e-06, 1.025813e-06, 1.04966e-06, 9.744175e-07, 1.012683e-06, 
    9.426047e-07, 9.629027e-07, 9.042791e-07, 9.331972e-07, 8.76836e-07, 
    8.53287e-07, 8.314386e-07, 8.062689e-07, 1.031732e-06, 1.040019e-06, 
    1.025206e-06, 1.004881e-06, 9.862108e-07, 9.61658e-07, 9.591648e-07, 
    9.54605e-07, 9.42848e-07, 9.330188e-07, 9.531632e-07, 9.305633e-07, 
    1.016804e-06, 9.711321e-07, 1.043158e-06, 1.021196e-06, 1.006074e-06, 
    1.012697e-06, 9.785517e-07, 9.705886e-07, 9.385669e-07, 9.550539e-07, 
    8.590662e-07, 9.008909e-07, 7.873845e-07, 8.183002e-07, 1.042921e-06, 
    1.031761e-06, 9.933816e-07, 1.011553e-06, 9.600313e-07, 9.47556e-07, 
    9.374776e-07, 9.2467e-07, 9.232944e-07, 9.157544e-07, 9.281263e-07, 
    9.162424e-07, 9.61606e-07, 9.411967e-07, 9.977348e-07, 9.838196e-07, 
    9.902099e-07, 9.972412e-07, 9.756202e-07, 9.528437e-07, 9.52364e-07, 
    9.451193e-07, 9.248486e-07, 9.598253e-07, 8.53736e-07, 9.184968e-07, 
    1.01966e-06, 9.984511e-07, 9.954448e-07, 1.003621e-06, 9.488029e-07, 
    9.68486e-07, 9.159383e-07, 9.299941e-07, 9.070221e-07, 9.184003e-07, 
    9.200803e-07, 9.348148e-07, 9.440473e-07, 9.675783e-07, 9.869408e-07, 
    1.002433e-06, 9.988206e-07, 9.818397e-07, 9.514602e-07, 9.231681e-07, 
    9.293279e-07, 9.087577e-07, 9.637214e-07, 9.404724e-07, 9.494229e-07, 
    9.261759e-07, 9.774984e-07, 9.33694e-07, 9.888561e-07, 9.839567e-07, 
    9.688788e-07, 9.389033e-07, 9.323418e-07, 9.253546e-07, 9.296638e-07, 
    9.50696e-07, 9.541662e-07, 9.692449e-07, 9.734272e-07, 9.850227e-07, 
    9.94673e-07, 9.85853e-07, 9.766321e-07, 9.506887e-07, 9.276096e-07, 
    9.027777e-07, 8.967548e-07, 8.682684e-07, 8.914164e-07, 8.533814e-07, 
    8.856558e-07, 8.301841e-07, 9.311925e-07, 8.86622e-07, 9.681969e-07, 
    9.592343e-07, 9.431262e-07, 9.067131e-07, 9.262846e-07, 9.034188e-07, 
    9.543027e-07, 9.812544e-07, 9.882941e-07, 1.001487e-06, 9.879934e-07, 
    9.890878e-07, 9.762539e-07, 9.803691e-07, 9.498335e-07, 9.661754e-07, 
    9.201215e-07, 9.035992e-07, 8.577745e-07, 8.302907e-07, 8.028001e-07, 
    7.908164e-07, 7.871881e-07, 7.856738e-07,
  8.152478e-08, 7.847274e-08, 7.906016e-08, 7.664195e-08, 7.797741e-08, 
    7.640269e-08, 8.089999e-08, 7.8353e-08, 7.997286e-08, 8.124712e-08, 
    7.2089e-08, 7.653526e-08, 6.765698e-08, 7.035664e-08, 6.370809e-08, 
    6.807226e-08, 6.285149e-08, 6.383163e-08, 6.091312e-08, 6.173988e-08, 
    5.810572e-08, 6.053406e-08, 5.628047e-08, 5.867973e-08, 5.829981e-08, 
    6.061526e-08, 7.562666e-08, 7.263286e-08, 7.580647e-08, 7.5374e-08, 
    7.556793e-08, 7.794954e-08, 7.9168e-08, 8.176147e-08, 8.128661e-08, 
    7.93839e-08, 7.518008e-08, 7.659044e-08, 7.306976e-08, 7.314807e-08, 
    6.935367e-08, 7.104786e-08, 6.486982e-08, 6.658777e-08, 6.170522e-08, 
    6.290967e-08, 6.176139e-08, 6.210812e-08, 6.175689e-08, 6.352971e-08, 
    6.2766e-08, 6.434129e-08, 7.072843e-08, 6.880927e-08, 7.463732e-08, 
    7.829355e-08, 8.078709e-08, 8.258751e-08, 8.23314e-08, 8.184453e-08, 
    7.937285e-08, 7.709457e-08, 7.53875e-08, 7.425962e-08, 7.315933e-08, 
    6.989389e-08, 6.820625e-08, 6.452592e-08, 6.518032e-08, 6.407453e-08, 
    6.303036e-08, 6.130269e-08, 6.158488e-08, 6.083152e-08, 6.410377e-08, 
    6.19161e-08, 6.555499e-08, 6.454582e-08, 7.286083e-08, 7.62083e-08, 
    7.766023e-08, 7.894698e-08, 8.21348e-08, 7.992443e-08, 8.079102e-08, 
    7.873969e-08, 7.745404e-08, 7.808821e-08, 7.422894e-08, 7.571393e-08, 
    6.810708e-08, 7.131815e-08, 6.315156e-08, 6.504567e-08, 6.270317e-08, 
    6.389136e-08, 6.18645e-08, 6.368668e-08, 6.055283e-08, 5.988434e-08, 
    6.03406e-08, 5.860102e-08, 6.37887e-08, 6.176128e-08, 7.810597e-08, 
    7.800229e-08, 7.752058e-08, 7.965271e-08, 7.978445e-08, 8.177445e-08, 
    8.000229e-08, 7.925526e-08, 7.738004e-08, 7.628451e-08, 7.525273e-08, 
    7.30167e-08, 7.057182e-08, 6.724555e-08, 6.492174e-08, 6.339446e-08, 
    6.432816e-08, 6.350335e-08, 6.442581e-08, 6.486129e-08, 6.013416e-08, 
    6.275884e-08, 5.884911e-08, 5.906109e-08, 6.081364e-08, 5.903718e-08, 
    7.792956e-08, 7.852705e-08, 8.06245e-08, 7.897997e-08, 8.199313e-08, 
    8.02972e-08, 7.933249e-08, 7.568242e-08, 7.489592e-08, 7.417108e-08, 
    7.275347e-08, 7.096048e-08, 6.788649e-08, 6.528538e-08, 6.297002e-08, 
    6.313779e-08, 6.307868e-08, 6.256837e-08, 6.383737e-08, 6.236168e-08, 
    6.211617e-08, 6.275929e-08, 5.908951e-08, 6.012279e-08, 5.90656e-08, 
    5.973685e-08, 7.833253e-08, 7.733059e-08, 7.787092e-08, 7.685684e-08, 
    7.757025e-08, 7.443084e-08, 7.350624e-08, 6.928124e-08, 7.099543e-08, 
    6.828071e-08, 7.071654e-08, 7.028071e-08, 6.819283e-08, 7.058354e-08, 
    6.54268e-08, 6.889395e-08, 6.254859e-08, 6.590862e-08, 6.234193e-08, 
    6.297991e-08, 6.192609e-08, 6.099226e-08, 5.983117e-08, 5.772773e-08, 
    5.821035e-08, 5.648051e-08, 7.585277e-08, 7.458207e-08, 7.469362e-08, 
    7.337785e-08, 7.241464e-08, 7.035612e-08, 6.713614e-08, 6.833528e-08, 
    6.614493e-08, 6.571086e-08, 6.904296e-08, 6.698387e-08, 7.373974e-08, 
    7.261868e-08, 7.328496e-08, 7.575188e-08, 6.805738e-08, 7.193777e-08, 
    6.488375e-08, 6.690312e-08, 6.112479e-08, 6.395452e-08, 5.847713e-08, 
    5.623491e-08, 5.41794e-08, 5.184157e-08, 7.38948e-08, 7.47514e-08, 
    7.322247e-08, 7.114107e-08, 6.924601e-08, 6.677872e-08, 6.652976e-08, 
    6.607523e-08, 6.490782e-08, 6.393691e-08, 6.593173e-08, 6.369508e-08, 
    7.235984e-08, 6.77274e-08, 7.507673e-08, 7.281039e-08, 7.126276e-08, 
    7.193918e-08, 6.847329e-08, 6.767286e-08, 6.448439e-08, 6.611993e-08, 
    5.678263e-08, 6.079593e-08, 5.010891e-08, 5.295503e-08, 7.505216e-08, 
    7.389786e-08, 6.997195e-08, 7.18222e-08, 6.661625e-08, 6.537452e-08, 
    6.437676e-08, 6.311589e-08, 6.298092e-08, 6.224283e-08, 6.345537e-08, 
    6.22905e-08, 6.677353e-08, 6.47444e-08, 7.041378e-08, 6.900448e-08, 
    6.965053e-08, 7.036363e-08, 6.817827e-08, 6.589995e-08, 6.58522e-08, 
    6.513285e-08, 6.313351e-08, 6.65957e-08, 5.627745e-08, 6.251104e-08, 
    7.265258e-08, 7.048661e-08, 7.018124e-08, 7.101264e-08, 6.54983e-08, 
    6.746201e-08, 6.226079e-08, 6.363907e-08, 6.139145e-08, 6.250152e-08, 
    6.266595e-08, 6.411396e-08, 6.502661e-08, 6.737105e-08, 6.93198e-08, 
    7.089169e-08, 7.052413e-08, 6.880468e-08, 6.576235e-08, 6.296855e-08, 
    6.357355e-08, 6.156036e-08, 6.698497e-08, 6.467276e-08, 6.555988e-08, 
    6.326373e-08, 6.836726e-08, 6.400354e-08, 6.95135e-08, 6.901831e-08, 
    6.750138e-08, 6.451765e-08, 6.387021e-08, 6.318309e-08, 6.360657e-08, 
    6.568638e-08, 6.603155e-08, 6.753807e-08, 6.795785e-08, 6.912595e-08, 
    7.010291e-08, 6.920985e-08, 6.828008e-08, 6.568564e-08, 6.340459e-08, 
    6.097898e-08, 6.039517e-08, 5.765821e-08, 5.987926e-08, 5.624389e-08, 
    5.932411e-08, 5.406218e-08, 6.375708e-08, 5.941707e-08, 6.743301e-08, 
    6.65367e-08, 6.493541e-08, 6.136142e-08, 6.32744e-08, 6.104124e-08, 
    6.604513e-08, 6.874568e-08, 6.945664e-08, 7.079539e-08, 6.942624e-08, 
    6.953695e-08, 6.824202e-08, 6.86564e-08, 6.560065e-08, 6.723053e-08, 
    6.266999e-08, 6.105876e-08, 5.666002e-08, 5.40721e-08, 5.152189e-08, 
    5.04224e-08, 5.009098e-08, 4.995285e-08,
  1.725263e-09, 1.63537e-09, 1.652568e-09, 1.582089e-09, 1.620906e-09, 
    1.575162e-09, 1.706753e-09, 1.631871e-09, 1.679388e-09, 1.71703e-09, 
    1.451727e-09, 1.578999e-09, 1.327853e-09, 1.402945e-09, 1.220101e-09, 
    1.339331e-09, 1.197062e-09, 1.223433e-09, 1.14538e-09, 1.167346e-09, 
    1.071661e-09, 1.135347e-09, 1.024467e-09, 1.086623e-09, 1.076713e-09, 
    1.137494e-09, 1.552751e-09, 1.467136e-09, 1.557936e-09, 1.545475e-09, 
    1.551059e-09, 1.620094e-09, 1.655731e-09, 1.732289e-09, 1.7182e-09, 
    1.662068e-09, 1.539896e-09, 1.580596e-09, 1.479545e-09, 1.481773e-09, 
    1.374914e-09, 1.422354e-09, 1.251538e-09, 1.29843e-09, 1.166423e-09, 
    1.198623e-09, 1.167919e-09, 1.177167e-09, 1.167799e-09, 1.215293e-09, 
    1.194769e-09, 1.237208e-09, 1.413375e-09, 1.359765e-09, 1.52431e-09, 
    1.630135e-09, 1.703414e-09, 1.756872e-09, 1.74924e-09, 1.734757e-09, 
    1.661743e-09, 1.595216e-09, 1.545863e-09, 1.513491e-09, 1.482093e-09, 
    1.389994e-09, 1.343039e-09, 1.242209e-09, 1.259978e-09, 1.229993e-09, 
    1.201862e-09, 1.155716e-09, 1.163219e-09, 1.143218e-09, 1.230783e-09, 
    1.172043e-09, 1.270183e-09, 1.242748e-09, 1.473609e-09, 1.56954e-09, 
    1.611664e-09, 1.649251e-09, 1.743388e-09, 1.677962e-09, 1.70353e-09, 
    1.643179e-09, 1.605663e-09, 1.624138e-09, 1.512613e-09, 1.555267e-09, 
    1.340294e-09, 1.429963e-09, 1.205118e-09, 1.256316e-09, 1.193085e-09, 
    1.225045e-09, 1.170667e-09, 1.219523e-09, 1.135844e-09, 1.118208e-09, 
    1.130236e-09, 1.084568e-09, 1.222275e-09, 1.167917e-09, 1.624657e-09, 
    1.621632e-09, 1.607598e-09, 1.669967e-09, 1.673842e-09, 1.732674e-09, 
    1.680254e-09, 1.658291e-09, 1.603511e-09, 1.571743e-09, 1.541985e-09, 
    1.478037e-09, 1.408979e-09, 1.31651e-09, 1.252948e-09, 1.211651e-09, 
    1.236852e-09, 1.214583e-09, 1.239497e-09, 1.251306e-09, 1.12479e-09, 
    1.194577e-09, 1.091049e-09, 1.096595e-09, 1.142745e-09, 1.095969e-09, 
    1.619511e-09, 1.636958e-09, 1.698609e-09, 1.650217e-09, 1.739173e-09, 
    1.688947e-09, 1.660558e-09, 1.554359e-09, 1.53173e-09, 1.510957e-09, 
    1.470558e-09, 1.419896e-09, 1.334192e-09, 1.262837e-09, 1.200242e-09, 
    1.204748e-09, 1.20316e-09, 1.189474e-09, 1.223588e-09, 1.183943e-09, 
    1.177382e-09, 1.194589e-09, 1.097339e-09, 1.12449e-09, 1.096713e-09, 
    1.114327e-09, 1.631272e-09, 1.602073e-09, 1.617802e-09, 1.588317e-09, 
    1.609044e-09, 1.518394e-09, 1.491974e-09, 1.372896e-09, 1.420879e-09, 
    1.345101e-09, 1.413041e-09, 1.400818e-09, 1.342668e-09, 1.409308e-09, 
    1.266689e-09, 1.362119e-09, 1.188944e-09, 1.279836e-09, 1.183414e-09, 
    1.200508e-09, 1.172309e-09, 1.147478e-09, 1.116809e-09, 1.061839e-09, 
    1.074383e-09, 1.02961e-09, 1.559272e-09, 1.522727e-09, 1.525925e-09, 
    1.488314e-09, 1.460947e-09, 1.40293e-09, 1.313497e-09, 1.346612e-09, 
    1.286297e-09, 1.274435e-09, 1.366262e-09, 1.309309e-09, 1.498633e-09, 
    1.466733e-09, 1.485669e-09, 1.556362e-09, 1.338918e-09, 1.44745e-09, 
    1.251916e-09, 1.307089e-09, 1.150993e-09, 1.226751e-09, 1.081335e-09, 
    1.023297e-09, 9.708782e-10, 9.122009e-10, 1.50306e-09, 1.527582e-09, 
    1.48389e-09, 1.424977e-09, 1.371914e-09, 1.303671e-09, 1.296839e-09, 
    1.28439e-09, 1.25257e-09, 1.226275e-09, 1.280467e-09, 1.219749e-09, 
    1.459395e-09, 1.329797e-09, 1.536924e-09, 1.472175e-09, 1.428403e-09, 
    1.447489e-09, 1.350438e-09, 1.328291e-09, 1.241084e-09, 1.285613e-09, 
    1.037393e-09, 1.142276e-09, 8.693735e-10, 9.400214e-10, 1.536218e-09, 
    1.503147e-09, 1.392175e-09, 1.444183e-09, 1.299211e-09, 1.265265e-09, 
    1.238168e-09, 1.20416e-09, 1.200535e-09, 1.180765e-09, 1.21329e-09, 
    1.18204e-09, 1.303529e-09, 1.248133e-09, 1.404546e-09, 1.365192e-09, 
    1.383194e-09, 1.403141e-09, 1.342264e-09, 1.279599e-09, 1.278294e-09, 
    1.258687e-09, 1.204635e-09, 1.298647e-09, 1.024391e-09, 1.187941e-09, 
    1.467694e-09, 1.406589e-09, 1.398032e-09, 1.421363e-09, 1.268637e-09, 
    1.322474e-09, 1.181246e-09, 1.218239e-09, 1.158075e-09, 1.187684e-09, 
    1.192087e-09, 1.231058e-09, 1.255798e-09, 1.319967e-09, 1.37397e-09, 
    1.417962e-09, 1.407641e-09, 1.359637e-09, 1.275841e-09, 1.200203e-09, 
    1.216474e-09, 1.162567e-09, 1.309339e-09, 1.24619e-09, 1.270316e-09, 
    1.208134e-09, 1.347499e-09, 1.228076e-09, 1.379371e-09, 1.365576e-09, 
    1.32356e-09, 1.241985e-09, 1.224474e-09, 1.205966e-09, 1.217363e-09, 
    1.273767e-09, 1.283196e-09, 1.324572e-09, 1.336165e-09, 1.368571e-09, 
    1.395839e-09, 1.370907e-09, 1.345083e-09, 1.273747e-09, 1.211924e-09, 
    1.147126e-09, 1.131677e-09, 1.060036e-09, 1.118075e-09, 1.023529e-09, 
    1.103489e-09, 9.679131e-10, 1.221422e-09, 1.105927e-09, 1.321674e-09, 
    1.297029e-09, 1.25332e-09, 1.157277e-09, 1.208421e-09, 1.148777e-09, 
    1.283567e-09, 1.357998e-09, 1.377785e-09, 1.415256e-09, 1.376937e-09, 
    1.380024e-09, 1.344029e-09, 1.355519e-09, 1.271428e-09, 1.316096e-09, 
    1.192196e-09, 1.149241e-09, 1.034232e-09, 9.681633e-10, 9.042557e-10, 
    8.770796e-10, 8.689331e-10, 8.655443e-10,
  1.149839e-11, 1.066681e-11, 1.08247e-11, 1.018137e-11, 1.053448e-11, 
    1.011867e-11, 1.132589e-11, 1.063476e-11, 1.107206e-11, 1.142158e-11, 
    9.018093e-12, 1.015339e-11, 7.946618e-12, 8.592058e-12, 7.043372e-12, 
    8.04444e-12, 6.853908e-12, 7.070883e-12, 6.433752e-12, 6.611493e-12, 
    5.846525e-12, 6.352989e-12, 5.478347e-12, 5.964531e-12, 5.886305e-12, 
    6.370252e-12, 9.916507e-12, 9.153734e-12, 9.963187e-12, 9.851083e-12, 
    9.901282e-12, 1.052705e-11, 1.085381e-11, 1.156403e-11, 1.143249e-11, 
    1.091216e-11, 9.800998e-12, 1.016785e-11, 9.263327e-12, 9.283035e-12, 
    8.349631e-12, 8.760933e-12, 7.304019e-12, 7.697228e-12, 6.604e-12, 
    6.866696e-12, 6.61615e-12, 6.691362e-12, 6.615175e-12, 7.003722e-12, 
    6.835121e-12, 7.184907e-12, 8.682709e-12, 8.21935e-12, 9.66142e-12, 
    1.061887e-11, 1.129484e-11, 1.179444e-11, 1.172279e-11, 1.158711e-11, 
    1.090917e-11, 1.030044e-11, 9.854569e-12, 9.564814e-12, 9.285872e-12, 
    8.479837e-12, 8.07611e-12, 7.22642e-12, 7.374401e-12, 7.125129e-12, 
    6.893273e-12, 6.517235e-12, 6.578007e-12, 6.416331e-12, 7.131664e-12, 
    6.649666e-12, 7.459732e-12, 7.230897e-12, 9.21086e-12, 1.006786e-11, 
    1.045014e-11, 1.07942e-11, 1.166792e-11, 1.105888e-11, 1.129593e-11, 
    1.073843e-11, 1.039545e-11, 1.056401e-11, 9.556985e-12, 9.939149e-12, 
    8.052661e-12, 8.827371e-12, 6.920008e-12, 7.343843e-12, 6.82133e-12, 
    7.084201e-12, 6.638478e-12, 7.038601e-12, 6.356977e-12, 6.215628e-12, 
    6.311948e-12, 5.94828e-12, 7.061315e-12, 6.61613e-12, 1.056875e-11, 
    1.05411e-11, 1.041308e-11, 1.098502e-11, 1.10208e-11, 1.156763e-11, 
    1.108008e-11, 1.087737e-11, 1.037586e-11, 1.008777e-11, 9.819744e-12, 
    9.249985e-12, 8.644475e-12, 7.850232e-12, 7.315766e-12, 6.973727e-12, 
    7.181957e-12, 6.997869e-12, 7.203895e-12, 7.302087e-12, 6.268286e-12, 
    6.83355e-12, 5.999552e-12, 6.043514e-12, 6.412516e-12, 6.038548e-12, 
    1.052173e-11, 1.068136e-11, 1.12502e-11, 1.080308e-11, 1.162844e-11, 
    1.116057e-11, 1.089825e-11, 9.930977e-12, 9.727806e-12, 9.542233e-12, 
    9.183911e-12, 8.739503e-12, 8.000606e-12, 7.398287e-12, 6.879978e-12, 
    6.916965e-12, 6.903924e-12, 6.79179e-12, 7.072161e-12, 6.746607e-12, 
    6.693116e-12, 6.833646e-12, 6.04942e-12, 6.265881e-12, 6.044451e-12, 
    6.18463e-12, 1.062927e-11, 1.036278e-11, 1.050612e-11, 1.023782e-11, 
    1.042625e-11, 9.608562e-12, 9.373431e-12, 8.332252e-12, 8.748071e-12, 
    8.093734e-12, 8.679802e-12, 8.573597e-12, 8.072944e-12, 8.647326e-12, 
    7.430497e-12, 8.239561e-12, 6.787461e-12, 7.540692e-12, 6.742295e-12, 
    6.882156e-12, 6.651827e-12, 6.450674e-12, 6.204443e-12, 5.76939e-12, 
    5.867948e-12, 5.518166e-12, 9.975222e-12, 9.647263e-12, 9.67585e-12, 
    9.340976e-12, 9.099177e-12, 8.591926e-12, 7.824687e-12, 8.106656e-12, 
    7.594986e-12, 7.495366e-12, 8.275157e-12, 7.789203e-12, 9.432562e-12, 
    9.150171e-12, 9.317537e-12, 9.949006e-12, 8.040919e-12, 8.980519e-12, 
    7.30717e-12, 7.770411e-12, 6.479054e-12, 7.098307e-12, 5.922753e-12, 
    5.469299e-12, 5.067949e-12, 4.628352e-12, 9.47192e-12, 9.690676e-12, 
    9.301778e-12, 8.783824e-12, 8.323792e-12, 7.741506e-12, 7.683801e-12, 
    7.578951e-12, 7.312613e-12, 7.094368e-12, 7.545988e-12, 7.040469e-12, 
    9.085525e-12, 7.963163e-12, 9.774349e-12, 9.198191e-12, 8.81374e-12, 
    8.980865e-12, 8.139395e-12, 7.950338e-12, 7.217073e-12, 7.589232e-12, 
    5.578567e-12, 6.408743e-12, 4.314222e-12, 4.835476e-12, 9.768017e-12, 
    9.472693e-12, 8.49871e-12, 8.951858e-12, 7.703825e-12, 7.418579e-12, 
    7.192873e-12, 6.912137e-12, 6.88238e-12, 6.720687e-12, 6.987225e-12, 
    6.731078e-12, 7.740301e-12, 7.275673e-12, 8.605957e-12, 8.265956e-12, 
    8.421058e-12, 8.593754e-12, 8.069482e-12, 7.538696e-12, 7.527737e-12, 
    7.363626e-12, 6.916049e-12, 7.699064e-12, 5.477764e-12, 6.779267e-12, 
    9.158643e-12, 8.623706e-12, 8.549436e-12, 8.752288e-12, 7.446795e-12, 
    7.90087e-12, 6.724601e-12, 7.028013e-12, 6.536321e-12, 6.777161e-12, 
    6.813169e-12, 7.133946e-12, 7.339521e-12, 7.879574e-12, 8.341498e-12, 
    8.722648e-12, 8.632838e-12, 8.218253e-12, 7.507155e-12, 6.879658e-12, 
    7.013459e-12, 6.572716e-12, 7.789455e-12, 7.259508e-12, 7.460856e-12, 
    6.944792e-12, 8.114238e-12, 7.109275e-12, 8.388053e-12, 8.269261e-12, 
    7.910098e-12, 7.224563e-12, 7.079484e-12, 6.926973e-12, 7.020789e-12, 
    7.489767e-12, 7.568912e-12, 7.9187e-12, 8.017426e-12, 8.295017e-12, 
    8.53043e-12, 8.31512e-12, 8.093583e-12, 7.489595e-12, 6.975975e-12, 
    6.447835e-12, 6.32351e-12, 5.755263e-12, 6.214566e-12, 5.471098e-12, 
    6.098293e-12, 5.045494e-12, 7.054284e-12, 6.117684e-12, 7.894076e-12, 
    7.685406e-12, 7.318866e-12, 6.52987e-12, 6.947152e-12, 6.461163e-12, 
    7.572031e-12, 8.204192e-12, 8.374374e-12, 8.699079e-12, 8.367063e-12, 
    8.393695e-12, 8.084564e-12, 8.182921e-12, 7.470165e-12, 7.846718e-12, 
    6.814056e-12, 6.464911e-12, 5.554016e-12, 5.047384e-12, 4.569636e-12, 
    4.370314e-12, 4.311022e-12, 4.28642e-12,
  1.443536e-14, 1.260027e-14, 1.294303e-14, 1.156368e-14, 1.231507e-14, 
    1.143176e-14, 1.404873e-14, 1.253102e-14, 1.348544e-14, 1.426282e-14, 
    9.192306e-15, 1.150475e-14, 7.162754e-15, 8.366476e-15, 5.582211e-15, 
    7.341379e-15, 5.267298e-15, 5.628429e-15, 4.591056e-15, 4.873329e-15, 
    3.700313e-15, 4.464687e-15, 3.176748e-15, 3.873967e-15, 3.758542e-15, 
    4.491599e-15, 1.100943e-14, 9.460209e-15, 1.110652e-14, 1.087379e-14, 
    1.097782e-14, 1.229914e-14, 1.300652e-14, 1.458327e-14, 1.42873e-14, 
    1.313406e-14, 1.077029e-14, 1.153519e-14, 9.678352e-15, 9.717746e-15, 
    7.907486e-15, 8.690933e-15, 6.025132e-15, 6.713758e-15, 4.861314e-15, 
    5.288358e-15, 4.8808e-15, 5.001998e-15, 4.879235e-15, 5.515804e-15, 
    5.2364e-15, 5.821347e-15, 8.540166e-15, 7.664201e-15, 1.048344e-14, 
    1.249674e-14, 1.397948e-14, 1.510595e-14, 1.494284e-14, 1.46354e-14, 
    1.312752e-14, 1.181548e-14, 1.0881e-14, 1.028628e-14, 9.723419e-15, 
    8.153016e-15, 7.399503e-15, 5.892115e-15, 6.146613e-15, 5.719946e-15, 
    5.332224e-15, 4.722931e-15, 4.819717e-15, 4.5637e-15, 5.731e-15, 
    4.934688e-15, 6.294945e-15, 5.899759e-15, 9.573743e-15, 1.132515e-14, 
    1.213434e-14, 1.28766e-14, 1.481828e-14, 1.345637e-14, 1.398189e-14, 
    1.27554e-14, 1.201756e-14, 1.237855e-14, 1.027035e-14, 1.105649e-14, 
    7.35645e-15, 8.819631e-15, 5.376473e-15, 6.09377e-15, 5.213757e-15, 
    5.650851e-15, 4.916678e-15, 5.5742e-15, 4.470902e-15, 4.252535e-15, 
    4.400933e-15, 3.849886e-15, 5.612338e-15, 4.880769e-15, 1.238874e-14, 
    1.23293e-14, 1.205516e-14, 1.329382e-14, 1.337249e-14, 1.459142e-14, 
    1.350313e-14, 1.305797e-14, 1.19758e-14, 1.136687e-14, 1.080899e-14, 
    9.651713e-15, 8.466776e-15, 6.988123e-15, 6.045351e-15, 5.465744e-15, 
    5.816327e-15, 5.506022e-15, 5.853679e-15, 6.021805e-15, 4.333449e-15, 
    5.23382e-15, 3.926032e-15, 3.99173e-15, 4.557717e-15, 3.984291e-15, 
    1.22877e-14, 1.263173e-14, 1.388006e-14, 1.289593e-14, 1.472886e-14, 
    1.368109e-14, 1.310363e-14, 1.10395e-14, 1.061958e-14, 1.024036e-14, 
    9.520105e-15, 8.649549e-15, 7.261159e-15, 6.188021e-15, 5.310264e-15, 
    5.371429e-15, 5.349837e-15, 5.165372e-15, 5.63058e-15, 5.091653e-15, 
    5.004838e-15, 5.233976e-15, 4.000585e-15, 4.32974e-15, 3.993135e-15, 
    4.205143e-15, 1.251916e-14, 1.194795e-14, 1.225421e-14, 1.168286e-14, 
    1.208328e-14, 1.037543e-14, 9.899072e-15, 7.874903e-15, 8.666089e-15, 
    7.431909e-15, 8.534577e-15, 8.331239e-15, 7.393691e-15, 8.472236e-15, 
    6.244004e-15, 7.701794e-15, 5.158293e-15, 6.43675e-15, 5.084636e-15, 
    5.31386e-15, 4.938165e-15, 4.617687e-15, 4.235412e-15, 3.588304e-15, 
    3.731628e-15, 3.232e-15, 1.113159e-14, 1.045448e-14, 1.051299e-14, 
    9.833847e-15, 9.352148e-15, 8.36622e-15, 6.94207e-15, 7.455695e-15, 
    6.532396e-15, 6.35723e-15, 7.768119e-15, 6.878267e-15, 1.001822e-14, 
    9.453126e-15, 9.786833e-15, 1.1077e-14, 7.334921e-15, 9.1185e-15, 
    6.030552e-15, 6.844548e-15, 4.662463e-15, 5.674638e-15, 3.81217e-15, 
    3.164244e-15, 2.627588e-15, 2.082997e-15, 1.009777e-14, 1.054337e-14, 
    9.755255e-15, 8.735216e-15, 7.859044e-15, 6.792795e-15, 6.689849e-15, 
    6.504099e-15, 6.03992e-15, 5.667988e-15, 6.446054e-15, 5.577333e-15, 
    9.325192e-15, 7.192861e-15, 1.071534e-14, 9.548512e-15, 8.793179e-15, 
    9.119169e-15, 7.516077e-15, 7.16951e-15, 5.876156e-15, 6.522235e-15, 
    3.316468e-15, 4.551804e-15, 1.72384e-15, 2.333719e-15, 1.07023e-14, 
    1.009933e-14, 8.188783e-15, 9.062328e-15, 6.725515e-15, 6.223265e-15, 
    5.834902e-15, 5.363434e-15, 5.31423e-15, 5.049523e-15, 5.488252e-15, 
    5.066398e-15, 6.790642e-15, 5.976426e-15, 8.393031e-15, 7.750958e-15, 
    8.041874e-15, 8.369711e-15, 7.387315e-15, 6.433237e-15, 6.41398e-15, 
    6.127965e-15, 5.369935e-15, 6.717029e-15, 3.175956e-15, 5.144923e-15, 
    9.469924e-15, 8.426995e-15, 8.285193e-15, 8.67423e-15, 6.272386e-15, 
    7.079692e-15, 5.055878e-15, 5.556451e-15, 4.753256e-15, 5.141464e-15, 
    5.200374e-15, 5.734862e-15, 6.08631e-15, 7.041135e-15, 7.892229e-15, 
    8.617037e-15, 8.44447e-15, 7.662163e-15, 6.377885e-15, 5.309739e-15, 
    5.532089e-15, 4.811264e-15, 6.878715e-15, 5.948714e-15, 6.296912e-15, 
    5.417599e-15, 7.469668e-15, 5.693167e-15, 7.979686e-15, 7.757118e-15, 
    7.09642e-15, 5.888946e-15, 5.642906e-15, 5.388021e-15, 5.544351e-15, 
    6.347433e-15, 6.486401e-15, 7.112022e-15, 7.291903e-15, 7.805207e-15, 
    8.249024e-15, 7.842806e-15, 7.43163e-15, 6.34713e-15, 5.469494e-15, 
    4.613217e-15, 4.418862e-15, 3.56793e-15, 4.250915e-15, 3.166741e-15, 
    4.074143e-15, 2.598655e-15, 5.600535e-15, 4.103435e-15, 7.06738e-15, 
    6.692705e-15, 6.050697e-15, 4.743006e-15, 5.421521e-15, 4.634223e-15, 
    6.491898e-15, 7.636055e-15, 7.953957e-15, 8.571647e-15, 7.940216e-15, 
    7.990306e-15, 7.415034e-15, 7.596599e-15, 6.313163e-15, 6.981777e-15, 
    5.201831e-15, 4.640134e-15, 3.282039e-15, 2.60108e-15, 2.01389e-15, 
    1.786039e-15, 1.720316e-15, 1.693328e-15,
  5.467353e-20, 4.78007e-20, 4.908537e-20, 4.391275e-20, 4.673143e-20, 
    4.34176e-20, 5.322654e-20, 4.75411e-20, 5.11174e-20, 5.402786e-20, 
    3.500043e-20, 4.369158e-20, 2.734916e-20, 3.189005e-20, 2.137153e-20, 
    2.802358e-20, 2.017821e-20, 2.15466e-20, 1.761264e-20, 1.868409e-20, 
    1.422577e-20, 1.71327e-20, 1.223033e-20, 1.488679e-20, 1.444746e-20, 
    1.723492e-20, 4.183204e-20, 3.600866e-20, 4.219662e-20, 4.132264e-20, 
    4.171334e-20, 4.667169e-20, 4.932328e-20, 5.522699e-20, 5.411946e-20, 
    4.980117e-20, 4.093389e-20, 4.380582e-20, 3.682934e-20, 3.697753e-20, 
    3.015963e-20, 3.311253e-20, 2.30486e-20, 2.565294e-20, 1.86385e-20, 
    2.025804e-20, 1.871244e-20, 1.917223e-20, 1.87065e-20, 2.111994e-20, 
    2.006108e-20, 2.227719e-20, 3.254455e-20, 2.924191e-20, 3.985618e-20, 
    4.741258e-20, 5.296729e-20, 5.718208e-20, 5.657203e-20, 5.542199e-20, 
    4.977664e-20, 4.485757e-20, 4.134972e-20, 3.91152e-20, 3.699886e-20, 
    3.108545e-20, 2.824299e-20, 2.254512e-20, 2.35083e-20, 2.189322e-20, 
    2.04243e-20, 1.811331e-20, 1.848065e-20, 1.750876e-20, 2.193508e-20, 
    1.891689e-20, 2.406945e-20, 2.257405e-20, 3.643582e-20, 4.301743e-20, 
    4.605368e-20, 4.883644e-20, 5.610616e-20, 5.100852e-20, 5.297633e-20, 
    4.838219e-20, 4.561564e-20, 4.696946e-20, 3.905534e-20, 4.200877e-20, 
    2.808047e-20, 3.359726e-20, 2.059199e-20, 2.330835e-20, 1.997525e-20, 
    2.163153e-20, 1.884857e-20, 2.134118e-20, 1.71563e-20, 1.632656e-20, 
    1.689049e-20, 1.479515e-20, 2.148565e-20, 1.871232e-20, 4.700769e-20, 
    4.678481e-20, 4.575669e-20, 5.039967e-20, 5.069437e-20, 5.525744e-20, 
    5.118366e-20, 4.951606e-20, 4.545902e-20, 4.317407e-20, 4.107925e-20, 
    3.672914e-20, 3.226802e-20, 2.66896e-20, 2.312512e-20, 2.093026e-20, 
    2.225819e-20, 2.108288e-20, 2.23996e-20, 2.303601e-20, 1.663408e-20, 
    2.005131e-20, 1.508491e-20, 1.533486e-20, 1.748603e-20, 1.530655e-20, 
    4.66288e-20, 4.791864e-20, 5.259509e-20, 4.890887e-20, 5.577163e-20, 
    5.185013e-20, 4.968716e-20, 4.194498e-20, 4.036769e-20, 3.894261e-20, 
    3.623402e-20, 3.295663e-20, 2.772072e-20, 2.366497e-20, 2.034107e-20, 
    2.057288e-20, 2.049105e-20, 1.97918e-20, 2.155475e-20, 1.951226e-20, 
    1.918301e-20, 2.00519e-20, 1.536854e-20, 1.661998e-20, 1.53402e-20, 
    1.614641e-20, 4.749666e-20, 4.535454e-20, 4.650323e-20, 4.435997e-20, 
    4.586219e-20, 3.945028e-20, 3.765948e-20, 3.003674e-20, 3.301894e-20, 
    2.836531e-20, 3.252349e-20, 3.175725e-20, 2.822105e-20, 3.228859e-20, 
    2.387676e-20, 2.938374e-20, 1.976496e-20, 2.460575e-20, 1.948565e-20, 
    2.03547e-20, 1.893008e-20, 1.771376e-20, 1.626148e-20, 1.379919e-20, 
    1.4345e-20, 1.24411e-20, 4.229076e-20, 3.974735e-20, 3.996719e-20, 
    3.741419e-20, 3.560202e-20, 3.188908e-20, 2.651563e-20, 2.845509e-20, 
    2.496739e-20, 2.430503e-20, 2.963395e-20, 2.627459e-20, 3.81075e-20, 
    3.5982e-20, 3.723738e-20, 4.208578e-20, 2.79992e-20, 3.47226e-20, 
    2.306912e-20, 2.614719e-20, 1.788376e-20, 2.172163e-20, 1.46516e-20, 
    1.218263e-20, 1.013288e-20, 8.047454e-21, 3.840658e-20, 4.008136e-20, 
    3.711861e-20, 3.327933e-20, 2.997693e-20, 2.595163e-20, 2.556258e-20, 
    2.48604e-20, 2.310457e-20, 2.169644e-20, 2.464093e-20, 2.135304e-20, 
    3.550058e-20, 2.746285e-20, 4.072747e-20, 3.63409e-20, 3.349764e-20, 
    3.472512e-20, 2.868298e-20, 2.737467e-20, 2.24847e-20, 2.492897e-20, 
    1.276322e-20, 1.746358e-20, 6.668523e-21, 9.008299e-21, 4.067846e-20, 
    3.841245e-20, 3.122028e-20, 3.451114e-20, 2.569738e-20, 2.37983e-20, 
    2.232851e-20, 2.054258e-20, 2.03561e-20, 1.935249e-20, 2.101554e-20, 
    1.941649e-20, 2.594349e-20, 2.286426e-20, 3.199012e-20, 2.956922e-20, 
    3.066641e-20, 3.190224e-20, 2.819698e-20, 2.459247e-20, 2.451964e-20, 
    2.343774e-20, 2.056722e-20, 2.566531e-20, 1.222731e-20, 1.971426e-20, 
    3.604522e-20, 3.211811e-20, 3.15837e-20, 3.304961e-20, 2.398412e-20, 
    2.703547e-20, 1.937659e-20, 2.127393e-20, 1.822842e-20, 1.970115e-20, 
    1.992451e-20, 2.194971e-20, 2.328012e-20, 2.688984e-20, 3.010209e-20, 
    3.283416e-20, 3.218397e-20, 2.923422e-20, 2.438314e-20, 2.033908e-20, 
    2.118163e-20, 1.844858e-20, 2.627628e-20, 2.275937e-20, 2.407689e-20, 
    2.074784e-20, 2.850782e-20, 2.17918e-20, 3.043191e-20, 2.959245e-20, 
    2.709865e-20, 2.253312e-20, 2.160144e-20, 2.063576e-20, 2.122809e-20, 
    2.426798e-20, 2.479349e-20, 2.715757e-20, 2.78368e-20, 2.977386e-20, 
    3.144737e-20, 2.991568e-20, 2.836426e-20, 2.426683e-20, 2.094447e-20, 
    1.769679e-20, 1.695861e-20, 1.372158e-20, 1.63204e-20, 1.219216e-20, 
    1.564831e-20, 1.002223e-20, 2.144094e-20, 1.575971e-20, 2.698897e-20, 
    2.557338e-20, 2.314536e-20, 1.818951e-20, 2.07627e-20, 1.777654e-20, 
    2.481427e-20, 2.913571e-20, 3.033488e-20, 3.266316e-20, 3.028307e-20, 
    3.047196e-20, 2.830161e-20, 2.898684e-20, 2.413836e-20, 2.666563e-20, 
    1.993003e-20, 1.779898e-20, 1.263194e-20, 1.003151e-20, 7.78237e-21, 
    6.907559e-21, 6.654977e-21, 6.551226e-21,
  4.403057e-26, 3.851807e-26, 3.954867e-26, 3.539844e-26, 3.76602e-26, 
    3.500107e-26, 4.287019e-26, 3.83098e-26, 4.117862e-26, 4.351281e-26, 
    2.824334e-26, 3.522095e-26, 2.209501e-26, 2.574466e-26, 1.728664e-26, 
    2.263722e-26, 1.632603e-26, 1.742755e-26, 1.425981e-26, 1.512287e-26, 
    1.152997e-26, 1.387313e-26, 9.920205e-27, 1.206298e-26, 1.170874e-26, 
    1.395549e-26, 3.372851e-26, 2.90531e-26, 3.402114e-26, 3.331963e-26, 
    3.363323e-26, 3.761227e-26, 3.973951e-26, 4.447437e-26, 4.358626e-26, 
    4.012286e-26, 3.300758e-26, 3.531263e-26, 2.971216e-26, 2.983116e-26, 
    2.435414e-26, 2.672683e-26, 1.86362e-26, 2.07311e-26, 1.508615e-26, 
    1.63903e-26, 1.51457e-26, 1.5516e-26, 1.514092e-26, 1.708415e-26, 
    1.623172e-26, 1.80155e-26, 2.627052e-26, 2.361655e-26, 3.214244e-26, 
    3.820669e-26, 4.266228e-26, 4.6042e-26, 4.555288e-26, 4.463074e-26, 
    4.010318e-26, 3.615664e-26, 3.334136e-26, 3.154757e-26, 2.984829e-26, 
    2.509814e-26, 2.28136e-26, 1.823109e-26, 1.900605e-26, 1.77065e-26, 
    1.652416e-26, 1.466313e-26, 1.495902e-26, 1.417612e-26, 1.774019e-26, 
    1.531037e-26, 1.945747e-26, 1.825437e-26, 2.939614e-26, 3.467992e-26, 
    3.711641e-26, 3.934897e-26, 4.517933e-26, 4.109129e-26, 4.266953e-26, 
    3.898457e-26, 3.676493e-26, 3.785117e-26, 3.149951e-26, 3.387036e-26, 
    2.268295e-26, 2.711624e-26, 1.665916e-26, 1.884518e-26, 1.616261e-26, 
    1.74959e-26, 1.525534e-26, 1.726222e-26, 1.389215e-26, 1.322354e-26, 
    1.367798e-26, 1.198909e-26, 1.737849e-26, 1.514561e-26, 3.788185e-26, 
    3.770302e-26, 3.687811e-26, 4.060293e-26, 4.083931e-26, 4.44988e-26, 
    4.123176e-26, 3.989416e-26, 3.663926e-26, 3.480562e-26, 3.312426e-26, 
    2.963169e-26, 2.604835e-26, 2.156471e-26, 1.869777e-26, 1.693147e-26, 
    1.80002e-26, 1.705432e-26, 1.8114e-26, 1.862607e-26, 1.347136e-26, 
    1.622385e-26, 1.222271e-26, 1.242421e-26, 1.415781e-26, 1.240139e-26, 
    3.757785e-26, 3.861269e-26, 4.236378e-26, 3.940708e-26, 4.49111e-26, 
    4.176631e-26, 4.00314e-26, 3.381916e-26, 3.255308e-26, 3.1409e-26, 
    2.923408e-26, 2.660159e-26, 2.239374e-26, 1.913208e-26, 1.645715e-26, 
    1.664377e-26, 1.65779e-26, 1.601491e-26, 1.74341e-26, 1.578982e-26, 
    1.552467e-26, 1.622433e-26, 1.245136e-26, 1.346e-26, 1.242851e-26, 
    1.307835e-26, 3.827415e-26, 3.655542e-26, 3.747711e-26, 3.575733e-26, 
    3.696276e-26, 3.181658e-26, 3.037876e-26, 2.425537e-26, 2.665164e-26, 
    2.291193e-26, 2.62536e-26, 2.563795e-26, 2.279596e-26, 2.606488e-26, 
    1.930246e-26, 2.373055e-26, 1.59933e-26, 1.988886e-26, 1.576839e-26, 
    1.646812e-26, 1.532099e-26, 1.434127e-26, 1.317109e-26, 1.118594e-26, 
    1.162612e-26, 1.009029e-26, 3.409669e-26, 3.205508e-26, 3.223156e-26, 
    3.01818e-26, 2.872652e-26, 2.574389e-26, 2.142483e-26, 2.29841e-26, 
    2.017974e-26, 1.964697e-26, 2.393166e-26, 2.1231e-26, 3.07385e-26, 
    2.903169e-26, 3.003982e-26, 3.393217e-26, 2.261762e-26, 2.802019e-26, 
    1.865271e-26, 2.112856e-26, 1.447822e-26, 1.756841e-26, 1.187335e-26, 
    9.881705e-27, 8.226696e-27, 6.541044e-27, 3.097863e-26, 3.232322e-26, 
    2.994445e-26, 2.686083e-26, 2.42073e-26, 2.09713e-26, 2.065843e-26, 
    2.009369e-26, 1.868123e-26, 1.754814e-26, 1.991716e-26, 1.727177e-26, 
    2.864505e-26, 2.218642e-26, 3.284188e-26, 2.931991e-26, 2.703621e-26, 
    2.802221e-26, 2.316728e-26, 2.211553e-26, 1.818248e-26, 2.014884e-26, 
    1.035021e-26, 1.413972e-26, 5.425151e-27, 7.317958e-27, 3.280254e-26, 
    3.098335e-26, 2.520649e-26, 2.785033e-26, 2.076683e-26, 1.923935e-26, 
    1.805679e-26, 1.661938e-26, 1.646925e-26, 1.566116e-26, 1.700012e-26, 
    1.571269e-26, 2.096475e-26, 1.848788e-26, 2.582507e-26, 2.387963e-26, 
    2.476141e-26, 2.575446e-26, 2.277661e-26, 1.987818e-26, 1.981961e-26, 
    1.894928e-26, 1.663921e-26, 2.074104e-26, 9.917763e-27, 1.595247e-26, 
    2.908245e-26, 2.592791e-26, 2.549851e-26, 2.667628e-26, 1.938883e-26, 
    2.184281e-26, 1.568057e-26, 1.72081e-26, 1.475585e-26, 1.594191e-26, 
    1.612176e-26, 1.775196e-26, 1.882247e-26, 2.172572e-26, 2.430789e-26, 
    2.650319e-26, 2.598082e-26, 2.361037e-26, 1.970981e-26, 1.645554e-26, 
    1.713381e-26, 1.493318e-26, 2.123236e-26, 1.840348e-26, 1.946346e-26, 
    1.678462e-26, 2.302649e-26, 1.762488e-26, 2.457296e-26, 2.38983e-26, 
    2.18936e-26, 1.822144e-26, 1.747168e-26, 1.669439e-26, 1.71712e-26, 
    1.961717e-26, 2.003987e-26, 2.194098e-26, 2.248706e-26, 2.40441e-26, 
    2.538896e-26, 2.415808e-26, 2.291108e-26, 1.961625e-26, 1.694291e-26, 
    1.43276e-26, 1.373286e-26, 1.112334e-26, 1.321858e-26, 9.889393e-27, 
    1.267688e-26, 8.137308e-27, 1.734251e-26, 1.276667e-26, 2.180542e-26, 
    2.066711e-26, 1.871404e-26, 1.472451e-26, 1.679659e-26, 1.439185e-26, 
    2.005659e-26, 2.353119e-26, 2.449498e-26, 2.636581e-26, 2.445334e-26, 
    2.460514e-26, 2.286072e-26, 2.341153e-26, 1.95129e-26, 2.154544e-26, 
    1.612621e-26, 1.440993e-26, 1.024428e-26, 8.144802e-27, 6.326617e-27, 
    5.618677e-27, 5.414182e-27, 5.330172e-27,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.00476365, 0.004763706, 0.004763696, 0.004763736, 0.004763716, 
    0.004763741, 0.004763664, 0.004763706, 0.004763681, 0.004763658, 
    0.004763797, 0.004763738, 0.004763922, 0.004763836, 0.004763969, 
    0.004763915, 0.004763979, 0.004763973, 0.004764003, 0.004763995, 
    0.004764016, 0.004764006, 0.004764031, 0.004764017, 0.004764018, 
    0.004764005, 0.004763756, 0.004763789, 0.004763753, 0.004763758, 
    0.004763757, 0.004763715, 0.004763689, 0.004763649, 0.004763657, 
    0.004763689, 0.004763761, 0.004763741, 0.004763799, 0.004763797, 
    0.00476385, 0.004763828, 0.004763961, 0.004763942, 0.004763996, 
    0.004763983, 0.004763994, 0.004763992, 0.004763994, 0.004763976, 
    0.004763984, 0.004763968, 0.004763831, 0.004763911, 0.004763771, 
    0.004763702, 0.004763665, 0.004763633, 0.004763637, 0.004763645, 
    0.004763689, 0.004763732, 0.004763762, 0.00476378, 0.004763797, 
    0.004763833, 0.004763915, 0.004763962, 0.004763959, 0.004763968, 
    0.004763982, 0.004763998, 0.004763996, 0.004764001, 0.004763971, 
    0.004763991, 0.004763956, 0.004763965, 0.004763785, 0.004763747, 
    0.004763715, 0.004763698, 0.00476364, 0.00476368, 0.004763664, 
    0.004763704, 0.004763726, 0.004763716, 0.00476378, 0.004763755, 
    0.004763917, 0.004763821, 0.00476398, 0.00476396, 0.004763986, 
    0.004763974, 0.004763992, 0.004763976, 0.004764005, 0.004764008, 
    0.004764006, 0.004764021, 0.004763974, 0.004763993, 0.004763715, 
    0.004763716, 0.004763726, 0.004763684, 0.004763682, 0.004763647, 
    0.004763681, 0.004763693, 0.004763728, 0.004763746, 0.004763762, 
    0.004763798, 0.004763831, 0.00476393, 0.004763961, 0.004763979, 
    0.004763969, 0.004763978, 0.004763968, 0.004763964, 0.004764006, 
    0.004763983, 0.004764019, 0.004764018, 0.004764001, 0.004764018, 
    0.004763718, 0.004763708, 0.004763668, 0.0047637, 0.004763644, 
    0.004763674, 0.004763689, 0.004763752, 0.004763769, 0.00476378, 
    0.004763803, 0.004763829, 0.004763923, 0.004763955, 0.004763984, 
    0.004763982, 0.004763982, 0.004763986, 0.004763973, 0.004763988, 
    0.004763989, 0.004763985, 0.004764018, 0.004764009, 0.004764018, 
    0.004764013, 0.004763712, 0.004763728, 0.004763719, 0.004763735, 
    0.004763722, 0.004763772, 0.004763785, 0.004763847, 0.004763827, 
    0.004763917, 0.004763832, 0.004763837, 0.004763911, 0.004763835, 
    0.00476395, 0.004763904, 0.004763986, 0.00476394, 0.004763989, 
    0.004763983, 0.004763994, 0.004764, 0.004764012, 0.004764024, 
    0.004764022, 0.004764033, 0.004763754, 0.004763771, 0.004763773, 
    0.004763793, 0.004763807, 0.004763838, 0.004763934, 0.00476392, 
    0.004763948, 0.004763952, 0.004763911, 0.004763934, 0.004763785, 
    0.004763799, 0.004763793, 0.004763753, 0.004763919, 0.004763809, 
    0.004763961, 0.004763938, 0.004763999, 0.004763968, 0.00476402, 
    0.004764026, 0.004764045, 0.004764043, 0.004763784, 0.004763772, 
    0.004763796, 0.004763822, 0.004763906, 0.004763938, 0.004763943, 
    0.004763948, 0.004763963, 0.004763973, 0.004763946, 0.004763976, 
    0.004763796, 0.004763925, 0.004763764, 0.004763796, 0.004763822, 
    0.004763814, 0.004763919, 0.004763929, 0.004763964, 0.004763949, 
    0.004764022, 0.004763997, 0.00476405, 0.004764043, 0.004763767, 
    0.004763786, 0.00476384, 0.004763816, 0.004763942, 0.004763956, 
    0.004763969, 0.004763979, 0.004763983, 0.004763989, 0.004763979, 
    0.00476399, 0.004763938, 0.004763964, 0.004763838, 0.00476391, 
    0.004763849, 0.004763839, 0.004763923, 0.004763945, 0.004763952, 
    0.004763957, 0.004763962, 0.004763943, 0.004764015, 0.00476397, 
    0.004763805, 0.00476383, 0.00476384, 0.00476383, 0.004763954, 0.00476393, 
    0.004763989, 0.004763976, 0.004763999, 0.004763987, 0.004763986, 
    0.004763971, 0.00476396, 0.004763931, 0.00476385, 0.004763831, 
    0.004763837, 0.004763911, 0.004763948, 0.004763981, 0.004763973, 
    0.004763997, 0.004763937, 0.004763962, 0.004763951, 0.004763979, 
    0.004763918, 0.004763955, 0.004763851, 0.004763911, 0.00476393, 
    0.00476396, 0.004763974, 0.004763979, 0.004763977, 0.00476395, 
    0.004763948, 0.004763931, 0.004763923, 0.004763911, 0.004763843, 
    0.004763908, 0.004763918, 0.004763952, 0.004763976, 0.004764, 
    0.004764007, 0.004764015, 0.004764002, 0.004764014, 0.004763993, 
    0.00476403, 0.004763965, 0.004764003, 0.004763932, 0.004763944, 
    0.004763957, 0.004763992, 0.004763979, 0.004763996, 0.004763948, 
    0.00476391, 0.004763851, 0.004763832, 0.004763851, 0.00476385, 
    0.004763922, 0.004763917, 0.004763953, 0.004763935, 0.004763984, 
    0.004763997, 0.00476403, 0.004764039, 0.004764051, 0.004764052, 
    0.004764053, 0.004764052,
  9.943882e-06, 9.95536e-06, 9.953137e-06, 9.962362e-06, 9.957258e-06, 
    9.963287e-06, 9.946224e-06, 9.955804e-06, 9.949698e-06, 9.944933e-06, 
    9.980171e-06, 9.962777e-06, 9.998363e-06, 9.987223e-06, 1.001506e-05, 
    9.996627e-06, 1.001877e-05, 1.001456e-05, 1.002729e-05, 1.002365e-05, 
    1.003983e-05, 1.002897e-05, 1.004824e-05, 1.003726e-05, 1.003897e-05, 
    1.002861e-05, 9.96631e-06, 9.978e-06, 9.96561e-06, 9.967281e-06, 
    9.966538e-06, 9.957354e-06, 9.952701e-06, 9.943023e-06, 9.944786e-06, 
    9.951904e-06, 9.968033e-06, 9.962583e-06, 9.976357e-06, 9.976048e-06, 
    9.991312e-06, 9.984436e-06, 1.001011e-05, 1.000286e-05, 1.00238e-05, 
    1.001854e-05, 1.002355e-05, 1.002203e-05, 1.002357e-05, 1.001585e-05, 
    1.001916e-05, 1.001237e-05, 9.98572e-06, 9.993621e-06, 9.970163e-06, 
    9.956002e-06, 9.94664e-06, 9.939962e-06, 9.940906e-06, 9.942701e-06, 
    9.951945e-06, 9.960642e-06, 9.967249e-06, 9.971659e-06, 9.976003e-06, 
    9.989051e-06, 9.996088e-06, 1.001156e-05, 1.00088e-05, 1.00135e-05, 
    1.001802e-05, 1.002556e-05, 1.002433e-05, 1.002764e-05, 1.001339e-05, 
    1.002286e-05, 1.000722e-05, 1.00115e-05, 9.977088e-06, 9.964058e-06, 
    9.958426e-06, 9.953561e-06, 9.94163e-06, 9.949868e-06, 9.946621e-06, 
    9.954363e-06, 9.959261e-06, 9.956843e-06, 9.971779e-06, 9.965976e-06, 
    9.996499e-06, 9.983331e-06, 1.001749e-05, 1.000937e-05, 1.001944e-05, 
    1.001431e-05, 1.002309e-05, 1.001519e-05, 1.002888e-05, 1.003184e-05, 
    1.002982e-05, 1.003763e-05, 1.001475e-05, 1.002354e-05, 9.956771e-06, 
    9.957164e-06, 9.959011e-06, 9.950889e-06, 9.950398e-06, 9.942969e-06, 
    9.949588e-06, 9.952396e-06, 9.959553e-06, 9.963762e-06, 9.967766e-06, 
    9.976558e-06, 9.986339e-06, 1.000009e-05, 1.000989e-05, 1.001645e-05, 
    1.001244e-05, 1.001598e-05, 1.001202e-05, 1.001016e-05, 1.003073e-05, 
    1.001918e-05, 1.003651e-05, 1.003556e-05, 1.002771e-05, 1.003566e-05, 
    9.957443e-06, 9.955173e-06, 9.947251e-06, 9.953452e-06, 9.94216e-06, 
    9.948472e-06, 9.952091e-06, 9.966076e-06, 9.969165e-06, 9.971998e-06, 
    9.97761e-06, 9.984788e-06, 9.99743e-06, 1.000834e-05, 1.001829e-05, 
    1.001756e-05, 1.001781e-05, 1.002002e-05, 1.001454e-05, 1.002092e-05, 
    1.002199e-05, 1.001919e-05, 1.003543e-05, 1.00308e-05, 1.003554e-05, 
    1.003252e-05, 9.955913e-06, 9.959736e-06, 9.957669e-06, 9.96155e-06, 
    9.958809e-06, 9.970956e-06, 9.97459e-06, 9.991583e-06, 9.984641e-06, 
    9.995794e-06, 9.985774e-06, 9.987531e-06, 9.996114e-06, 9.986318e-06, 
    1.000772e-05, 9.993244e-06, 1.002011e-05, 1.000566e-05, 1.002101e-05, 
    1.001824e-05, 1.002283e-05, 1.002693e-05, 1.00321e-05, 1.004158e-05, 
    1.003939e-05, 1.004733e-05, 9.965437e-06, 9.970376e-06, 9.969958e-06, 
    9.975133e-06, 9.978951e-06, 9.987238e-06, 1.000056e-05, 9.995591e-06, 
    1.000472e-05, 1.000655e-05, 9.992684e-06, 1.000118e-05, 9.97369e-06, 
    9.978113e-06, 9.975493e-06, 9.965816e-06, 9.996712e-06, 9.980833e-06, 
    1.001005e-05, 1.000154e-05, 1.002635e-05, 1.001401e-05, 1.003818e-05, 
    1.004843e-05, 1.005812e-05, 1.006933e-05, 9.973087e-06, 9.969733e-06, 
    9.975753e-06, 9.984034e-06, 9.99184e-06, 1.000205e-05, 1.000311e-05, 
    1.000501e-05, 1.000996e-05, 1.001411e-05, 1.000559e-05, 1.001515e-05, 
    9.979101e-06, 9.998088e-06, 9.968448e-06, 9.977345e-06, 9.983555e-06, 
    9.98085e-06, 9.995028e-06, 9.998336e-06, 1.001174e-05, 1.000483e-05, 
    1.004588e-05, 1.002777e-05, 1.00779e-05, 1.006394e-05, 9.968556e-06, 
    9.973084e-06, 9.988779e-06, 9.981321e-06, 1.000274e-05, 1.000797e-05, 
    1.001223e-05, 1.001764e-05, 1.001823e-05, 1.002144e-05, 1.001619e-05, 
    1.002124e-05, 1.000207e-05, 1.001065e-05, 9.987009e-06, 9.99283e-06, 
    9.990114e-06, 9.987212e-06, 9.996244e-06, 1.000572e-05, 1.000596e-05, 
    1.000899e-05, 1.001746e-05, 1.000283e-05, 1.004816e-05, 1.002018e-05, 
    9.978015e-06, 9.986672e-06, 9.987943e-06, 9.984586e-06, 1.000744e-05, 
    9.999204e-06, 1.002136e-05, 1.001539e-05, 1.002518e-05, 1.002032e-05, 
    1.00196e-05, 1.001335e-05, 1.000945e-05, 9.999577e-06, 9.99145e-06, 
    9.985077e-06, 9.986562e-06, 9.993645e-06, 1.000631e-05, 1.001828e-05, 
    1.001565e-05, 1.002444e-05, 1.00012e-05, 1.001094e-05, 1.000717e-05, 
    1.001701e-05, 9.995453e-06, 1.001373e-05, 9.990674e-06, 9.992784e-06, 
    9.99904e-06, 1.001158e-05, 1.00144e-05, 1.001735e-05, 1.001553e-05, 
    1.000664e-05, 1.000519e-05, 9.998896e-06, 9.997141e-06, 9.992345e-06, 
    9.988272e-06, 9.991993e-06, 9.995804e-06, 1.000665e-05, 1.001639e-05, 
    1.002699e-05, 1.002959e-05, 1.004185e-05, 1.003183e-05, 1.004831e-05, 
    1.003424e-05, 1.005859e-05, 1.001483e-05, 1.003389e-05, 9.999335e-06, 
    1.000308e-05, 1.000981e-05, 1.002527e-05, 1.001696e-05, 1.002669e-05, 
    1.000514e-05, 9.993872e-06, 9.990904e-06, 9.985459e-06, 9.991028e-06, 
    9.990576e-06, 9.995983e-06, 9.994274e-06, 1.000701e-05, 1.000018e-05, 
    1.001957e-05, 1.002662e-05, 1.004649e-05, 1.00586e-05, 1.007094e-05, 
    1.007635e-05, 1.0078e-05, 1.007869e-05,
  2.187819e-10, 2.192561e-10, 2.191641e-10, 2.19546e-10, 2.193345e-10, 
    2.195843e-10, 2.188785e-10, 2.192745e-10, 2.190219e-10, 2.188252e-10, 
    2.202857e-10, 2.195632e-10, 2.210414e-10, 2.205788e-10, 2.217398e-10, 
    2.20969e-10, 2.218954e-10, 2.217186e-10, 2.222531e-10, 2.221e-10, 
    2.227814e-10, 2.223237e-10, 2.23136e-10, 2.226726e-10, 2.227447e-10, 
    2.223084e-10, 2.197095e-10, 2.201954e-10, 2.196805e-10, 2.197499e-10, 
    2.19719e-10, 2.193386e-10, 2.191462e-10, 2.187463e-10, 2.188191e-10, 
    2.191132e-10, 2.197811e-10, 2.19555e-10, 2.201266e-10, 2.201137e-10, 
    2.207492e-10, 2.204626e-10, 2.215325e-10, 2.212291e-10, 2.221064e-10, 
    2.218857e-10, 2.220959e-10, 2.220323e-10, 2.220967e-10, 2.21773e-10, 
    2.219117e-10, 2.216271e-10, 2.205161e-10, 2.208434e-10, 2.198694e-10, 
    2.192829e-10, 2.188957e-10, 2.186201e-10, 2.18659e-10, 2.187331e-10, 
    2.191149e-10, 2.194746e-10, 2.197484e-10, 2.199314e-10, 2.201118e-10, 
    2.206553e-10, 2.209464e-10, 2.215933e-10, 2.214774e-10, 2.216744e-10, 
    2.218638e-10, 2.221805e-10, 2.221285e-10, 2.222678e-10, 2.216698e-10, 
    2.22067e-10, 2.214112e-10, 2.215905e-10, 2.201576e-10, 2.196162e-10, 
    2.193832e-10, 2.191817e-10, 2.186889e-10, 2.19029e-10, 2.188949e-10, 
    2.192147e-10, 2.194174e-10, 2.193173e-10, 2.199364e-10, 2.196956e-10, 
    2.209636e-10, 2.204168e-10, 2.218417e-10, 2.215013e-10, 2.219234e-10, 
    2.217082e-10, 2.220766e-10, 2.217451e-10, 2.2232e-10, 2.224447e-10, 
    2.223594e-10, 2.226883e-10, 2.217266e-10, 2.220956e-10, 2.193144e-10, 
    2.193307e-10, 2.19407e-10, 2.190713e-10, 2.190509e-10, 2.187441e-10, 
    2.190174e-10, 2.191335e-10, 2.194295e-10, 2.196039e-10, 2.197699e-10, 
    2.20135e-10, 2.20542e-10, 2.211134e-10, 2.215233e-10, 2.217979e-10, 
    2.216298e-10, 2.217782e-10, 2.216121e-10, 2.215344e-10, 2.223978e-10, 
    2.219128e-10, 2.22641e-10, 2.226008e-10, 2.22271e-10, 2.226054e-10, 
    2.193422e-10, 2.192482e-10, 2.189209e-10, 2.191771e-10, 2.187108e-10, 
    2.189714e-10, 2.19121e-10, 2.196999e-10, 2.198279e-10, 2.199455e-10, 
    2.201786e-10, 2.204773e-10, 2.210023e-10, 2.214583e-10, 2.218749e-10, 
    2.218445e-10, 2.218552e-10, 2.219479e-10, 2.217177e-10, 2.219857e-10, 
    2.220303e-10, 2.219131e-10, 2.225954e-10, 2.224006e-10, 2.226e-10, 
    2.224732e-10, 2.192788e-10, 2.194371e-10, 2.193515e-10, 2.195123e-10, 
    2.193988e-10, 2.199024e-10, 2.200534e-10, 2.207606e-10, 2.204712e-10, 
    2.20934e-10, 2.205184e-10, 2.205916e-10, 2.209477e-10, 2.20541e-10, 
    2.214325e-10, 2.208278e-10, 2.219515e-10, 2.213465e-10, 2.219893e-10, 
    2.218731e-10, 2.220658e-10, 2.22238e-10, 2.224553e-10, 2.22855e-10, 
    2.227626e-10, 2.230974e-10, 2.196733e-10, 2.198783e-10, 2.198608e-10, 
    2.200757e-10, 2.202345e-10, 2.205793e-10, 2.211329e-10, 2.209254e-10, 
    2.213069e-10, 2.213833e-10, 2.208041e-10, 2.211591e-10, 2.200159e-10, 
    2.201997e-10, 2.200907e-10, 2.196891e-10, 2.209724e-10, 2.203129e-10, 
    2.2153e-10, 2.211737e-10, 2.222134e-10, 2.216958e-10, 2.227116e-10, 
    2.23144e-10, 2.235537e-10, 2.240289e-10, 2.199908e-10, 2.198515e-10, 
    2.201014e-10, 2.204461e-10, 2.20769e-10, 2.211953e-10, 2.212393e-10, 
    2.21319e-10, 2.215261e-10, 2.216999e-10, 2.213435e-10, 2.217436e-10, 
    2.202412e-10, 2.210298e-10, 2.197982e-10, 2.201679e-10, 2.204261e-10, 
    2.203134e-10, 2.209019e-10, 2.2104e-10, 2.216009e-10, 2.213114e-10, 
    2.230367e-10, 2.222735e-10, 2.243928e-10, 2.238005e-10, 2.198026e-10, 
    2.199906e-10, 2.206436e-10, 2.20333e-10, 2.212241e-10, 2.214428e-10, 
    2.21621e-10, 2.218479e-10, 2.218728e-10, 2.220073e-10, 2.217869e-10, 
    2.219988e-10, 2.211962e-10, 2.21555e-10, 2.205698e-10, 2.208103e-10, 
    2.206991e-10, 2.205782e-10, 2.209526e-10, 2.21349e-10, 2.213585e-10, 
    2.214854e-10, 2.218411e-10, 2.212277e-10, 2.231333e-10, 2.21955e-10, 
    2.201954e-10, 2.20556e-10, 2.206087e-10, 2.204688e-10, 2.214208e-10, 
    2.210763e-10, 2.220042e-10, 2.217537e-10, 2.221643e-10, 2.219602e-10, 
    2.219301e-10, 2.216681e-10, 2.215047e-10, 2.210919e-10, 2.207549e-10, 
    2.204892e-10, 2.205511e-10, 2.208443e-10, 2.213735e-10, 2.218746e-10, 
    2.217647e-10, 2.221331e-10, 2.211596e-10, 2.215674e-10, 2.214094e-10, 
    2.218214e-10, 2.209197e-10, 2.216845e-10, 2.207225e-10, 2.208083e-10, 
    2.210695e-10, 2.215943e-10, 2.217119e-10, 2.218357e-10, 2.217595e-10, 
    2.213871e-10, 2.213265e-10, 2.210634e-10, 2.209902e-10, 2.2079e-10, 
    2.206223e-10, 2.207754e-10, 2.209344e-10, 2.213877e-10, 2.217955e-10, 
    2.222403e-10, 2.223496e-10, 2.228666e-10, 2.224443e-10, 2.231397e-10, 
    2.225464e-10, 2.235742e-10, 2.217303e-10, 2.22531e-10, 2.210817e-10, 
    2.212381e-10, 2.2152e-10, 2.221684e-10, 2.218195e-10, 2.222281e-10, 
    2.213242e-10, 2.208539e-10, 2.207321e-10, 2.205052e-10, 2.207372e-10, 
    2.207184e-10, 2.209417e-10, 2.208704e-10, 2.214027e-10, 2.211169e-10, 
    2.219291e-10, 2.222251e-10, 2.23062e-10, 2.235741e-10, 2.240968e-10, 
    2.24327e-10, 2.243971e-10, 2.244264e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  2.496702, 2.473692, 2.478171, 2.459571, 2.469895, 2.457708, 2.492044, 
    2.472776, 2.485082, 2.494635, 2.423349, 2.458741, 2.386433, 2.409123, 
    2.352012, 2.389967, 2.344339, 2.353112, 2.326687, 2.334265, 2.300374, 
    2.323187, 2.282759, 2.305829, 2.302222, 2.323938, 2.451633, 2.427763, 
    2.453045, 2.449646, 2.451172, 2.469681, 2.478991, 2.49846, 2.49493, 
    2.480629, 2.448117, 2.45917, 2.43129, 2.431921, 2.400769, 2.414829, 
    2.362297, 2.377262, 2.333949, 2.344862, 2.334462, 2.337617, 2.33442, 
    2.35042, 2.343568, 2.357635, 2.412197, 2.396198, 2.443823, 2.472321, 
    2.491199, 2.504566, 2.502677, 2.499076, 2.480546, 2.463085, 2.449752, 
    2.440821, 2.432011, 2.405281, 2.391103, 2.359267, 2.365023, 2.355271, 
    2.345947, 2.330267, 2.33285, 2.325935, 2.35553, 2.335871, 2.3683, 
    2.359442, 2.429606, 2.45619, 2.467456, 2.47731, 2.501225, 2.484717, 
    2.491229, 2.47573, 2.465865, 2.470746, 2.440576, 2.452319, 2.390262, 
    2.41705, 2.347035, 2.363842, 2.343002, 2.353643, 2.335402, 2.35182, 
    2.32336, 2.31715, 2.321394, 2.305083, 2.35273, 2.334461, 2.470882, 
    2.470086, 2.466378, 2.482665, 2.48366, 2.498556, 2.485304, 2.479653, 
    2.465293, 2.456785, 2.44869, 2.430862, 2.410904, 2.382917, 2.362754, 
    2.349211, 2.357518, 2.350184, 2.358382, 2.362222, 2.319477, 2.343504, 
    2.307431, 2.309431, 2.32577, 2.309205, 2.469527, 2.474107, 2.489981, 
    2.477561, 2.500177, 2.487525, 2.480239, 2.452072, 2.445872, 2.440115, 
    2.428737, 2.41411, 2.388388, 2.365944, 2.345405, 2.346911, 2.346381, 
    2.341785, 2.353163, 2.339916, 2.33769, 2.343508, 2.309699, 2.319371, 
    2.309473, 2.315773, 2.472619, 2.464911, 2.469077, 2.461241, 2.466762, 
    2.442183, 2.4348, 2.400163, 2.414398, 2.391734, 2.412099, 2.408494, 
    2.39099, 2.411, 2.367181, 2.396911, 2.341607, 2.371381, 2.339737, 
    2.345494, 2.335962, 2.327415, 2.316654, 2.296759, 2.30137, 2.284709, 
    2.453408, 2.443385, 2.444269, 2.433769, 2.425994, 2.409118, 2.381979, 
    2.392195, 2.373432, 2.369659, 2.398163, 2.380672, 2.436671, 2.427647, 
    2.433022, 2.452617, 2.38984, 2.422117, 2.36242, 2.379978, 2.328635, 
    2.354205, 2.303907, 2.282314, 2.261953, 2.238092, 2.437911, 2.444727, 
    2.432519, 2.415596, 2.399867, 2.378908, 2.376761, 2.372827, 2.362631, 
    2.354048, 2.371582, 2.351895, 2.42555, 2.387033, 2.447301, 2.429198, 
    2.416595, 2.422128, 2.393363, 2.386568, 2.3589, 2.373215, 2.287647, 
    2.325607, 2.21989, 2.249554, 2.447107, 2.437935, 2.405929, 2.421174, 
    2.377507, 2.366724, 2.357948, 2.346715, 2.345503, 2.338839, 2.349755, 
    2.339272, 2.378863, 2.361193, 2.409596, 2.39784, 2.403251, 2.409181, 
    2.390865, 2.371305, 2.37089, 2.364607, 2.346875, 2.37733, 2.282731, 
    2.341269, 2.427921, 2.4102, 2.407668, 2.414539, 2.367805, 2.384768, 
    2.339002, 2.351396, 2.331081, 2.341181, 2.342666, 2.35562, 2.363675, 
    2.383991, 2.400486, 2.413543, 2.410509, 2.396159, 2.370108, 2.345392, 
    2.350811, 2.332626, 2.380681, 2.360562, 2.368343, 2.348041, 2.392466, 
    2.354642, 2.402106, 2.397956, 2.385105, 2.359194, 2.353455, 2.347318, 
    2.351106, 2.369446, 2.372448, 2.385418, 2.388994, 2.39886, 2.407018, 
    2.399564, 2.391728, 2.36944, 2.349302, 2.327293, 2.3219, 2.296093, 
    2.317103, 2.282403, 2.311908, 2.260776, 2.352449, 2.312779, 2.384521, 
    2.376821, 2.362874, 2.330806, 2.348136, 2.327867, 2.372566, 2.395662, 
    2.401631, 2.41275, 2.401376, 2.402302, 2.391406, 2.394909, 2.368699, 
    2.382788, 2.342703, 2.328028, 2.286456, 2.260875, 2.234767, 2.223217, 
    2.219699, 2.218228,
  1.658923, 1.637599, 1.641748, 1.624528, 1.634084, 1.622804, 1.654604, 
    1.636751, 1.648152, 1.657007, 1.591043, 1.62376, 1.556995, 1.577915, 
    1.525317, 1.56025, 1.518266, 1.526329, 1.502058, 1.509014, 1.47793, 
    1.498846, 1.461804, 1.482929, 1.479624, 1.499535, 1.617185, 1.595119, 
    1.61849, 1.615346, 1.616758, 1.633886, 1.642507, 1.660553, 1.65728, 
    1.644025, 1.613932, 1.624157, 1.59838, 1.598963, 1.57021, 1.583181, 
    1.534777, 1.548549, 1.508724, 1.518747, 1.509194, 1.512092, 1.509157, 
    1.523855, 1.517559, 1.530488, 1.580752, 1.565995, 1.609962, 1.636329, 
    1.653821, 1.666216, 1.664465, 1.661124, 1.643948, 1.62778, 1.615445, 
    1.607187, 1.599046, 1.574368, 1.561298, 1.531989, 1.537285, 1.528314, 
    1.519744, 1.505344, 1.507715, 1.501367, 1.528553, 1.510489, 1.5403, 
    1.532151, 1.596821, 1.6214, 1.631824, 1.640951, 1.663118, 1.647813, 
    1.653848, 1.639488, 1.630353, 1.634872, 1.606961, 1.617819, 1.560523, 
    1.585229, 1.520744, 1.536198, 1.517038, 1.526818, 1.510057, 1.525143, 
    1.499005, 1.493308, 1.497201, 1.482246, 1.525978, 1.509193, 1.634998, 
    1.634261, 1.630829, 1.645911, 1.646834, 1.660643, 1.648357, 1.643121, 
    1.629824, 1.621951, 1.614463, 1.597985, 1.579558, 1.553756, 1.535196, 
    1.522744, 1.530381, 1.523639, 1.531176, 1.534708, 1.495442, 1.517499, 
    1.484397, 1.486231, 1.501216, 1.486024, 1.633744, 1.637984, 1.652692, 
    1.641183, 1.662145, 1.650415, 1.643664, 1.617589, 1.611857, 1.606535, 
    1.596022, 1.582517, 1.558796, 1.538131, 1.519246, 1.520631, 1.520143, 
    1.515921, 1.526376, 1.514204, 1.512159, 1.517503, 1.486476, 1.495345, 
    1.48627, 1.492045, 1.636606, 1.62947, 1.633327, 1.626074, 1.631183, 
    1.608446, 1.601622, 1.56965, 1.582782, 1.56188, 1.580661, 1.577334, 
    1.561193, 1.579648, 1.539269, 1.566651, 1.515757, 1.543133, 1.51404, 
    1.519328, 1.510572, 1.502726, 1.492853, 1.47462, 1.478844, 1.463589, 
    1.618826, 1.609557, 1.610375, 1.60067, 1.593488, 1.577911, 1.552893, 
    1.562306, 1.545023, 1.541551, 1.567807, 1.551689, 1.603351, 1.595014, 
    1.59998, 1.618094, 1.560134, 1.589907, 1.534889, 1.55105, 1.503845, 
    1.527334, 1.481168, 1.461396, 1.442784, 1.421004, 1.604497, 1.610799, 
    1.599516, 1.583887, 1.569378, 1.550064, 1.548088, 1.544466, 1.535084, 
    1.527191, 1.543319, 1.525212, 1.593076, 1.557548, 1.613178, 1.596446, 
    1.58481, 1.589918, 1.563382, 1.557121, 1.531651, 1.544824, 1.466276, 
    1.501065, 1.404418, 1.431461, 1.612999, 1.60452, 1.574968, 1.589037, 
    1.548775, 1.538849, 1.530777, 1.52045, 1.519336, 1.513215, 1.523245, 
    1.513612, 1.550023, 1.533761, 1.578352, 1.567509, 1.572499, 1.577969, 
    1.56108, 1.543065, 1.542683, 1.536901, 1.520593, 1.548612, 1.461775, 
    1.515443, 1.595268, 1.578907, 1.576573, 1.582913, 1.539844, 1.555462, 
    1.513364, 1.524752, 1.506091, 1.515366, 1.51673, 1.528636, 1.536044, 
    1.554746, 1.569948, 1.581994, 1.579194, 1.565959, 1.541963, 1.519234, 
    1.524215, 1.507509, 1.551698, 1.53318, 1.540339, 1.521668, 1.562555, 
    1.527733, 1.571443, 1.567616, 1.555772, 1.531921, 1.526645, 1.521004, 
    1.524486, 1.541354, 1.544117, 1.556061, 1.559356, 1.56845, 1.575973, 
    1.569098, 1.561875, 1.541348, 1.522827, 1.502614, 1.497666, 1.474009, 
    1.493263, 1.461475, 1.488497, 1.441706, 1.525718, 1.489298, 1.555234, 
    1.548143, 1.535306, 1.505837, 1.521756, 1.503139, 1.544226, 1.5655, 
    1.571005, 1.581262, 1.57077, 1.571624, 1.561578, 1.564807, 1.540666, 
    1.553638, 1.516763, 1.503287, 1.465187, 1.441798, 1.417974, 1.407449, 
    1.404245, 1.402905,
  0.6537162, 0.642145, 0.6443916, 0.6350822, 0.6402435, 0.6341522, 0.6513676, 
    0.6416858, 0.6478635, 0.6526738, 0.6170963, 0.6346678, 0.598967, 
    0.6100869, 0.5822451, 0.6006933, 0.5785421, 0.5827771, 0.5700572, 
    0.5736944, 0.5574961, 0.5683804, 0.5491477, 0.5600916, 0.5583754, 
    0.5687401, 0.6311247, 0.6192775, 0.6318278, 0.6301351, 0.6308949, 
    0.6401362, 0.6448027, 0.6546035, 0.6528223, 0.6456255, 0.6293744, 
    0.6348823, 0.6210241, 0.6213363, 0.6059841, 0.6128955, 0.5872235, 
    0.5944947, 0.5735425, 0.5787947, 0.5737886, 0.5753057, 0.5737689, 
    0.5814765, 0.5781711, 0.5849649, 0.6115994, 0.6037431, 0.6272394, 
    0.6414575, 0.6509421, 0.6576882, 0.6567336, 0.6549143, 0.6455835, 
    0.6368372, 0.6301883, 0.6257487, 0.6213812, 0.6081976, 0.6012492, 
    0.5857549, 0.5885456, 0.5838209, 0.5793179, 0.5717744, 0.5730146, 
    0.5696966, 0.5839466, 0.574466, 0.5901363, 0.5858402, 0.6201891, 
    0.6333957, 0.6390218, 0.6439594, 0.6559998, 0.6476797, 0.6509569, 
    0.6431672, 0.6382268, 0.6406695, 0.6256274, 0.6314662, 0.6008379, 
    0.6139894, 0.5798427, 0.5879727, 0.5778982, 0.5830341, 0.5742402, 
    0.5821533, 0.5684634, 0.5654924, 0.5675222, 0.5597367, 0.5825925, 
    0.5737881, 0.6407377, 0.6403391, 0.6384836, 0.646648, 0.6471485, 
    0.6546521, 0.6479751, 0.6451356, 0.6379411, 0.6336924, 0.6296597, 
    0.6208122, 0.6109627, 0.5972508, 0.5874448, 0.5808929, 0.5849088, 
    0.5813629, 0.5853269, 0.5871872, 0.5666048, 0.57814, 0.5608549, 
    0.5618082, 0.5696176, 0.5617008, 0.6400594, 0.6423533, 0.6503288, 
    0.6440855, 0.6554703, 0.6490919, 0.6454297, 0.6313427, 0.6282579, 
    0.6253985, 0.6197608, 0.6125413, 0.5999219, 0.588992, 0.5790564, 
    0.5797831, 0.5795272, 0.5773121, 0.5828019, 0.5764121, 0.5753407, 
    0.578142, 0.5619358, 0.5665544, 0.5618284, 0.5648345, 0.6416076, 0.63775, 
    0.6398338, 0.6359162, 0.6386752, 0.6264248, 0.6227618, 0.6056863, 
    0.6126829, 0.6015579, 0.6115512, 0.6097775, 0.6011933, 0.6110106, 
    0.5895923, 0.6040921, 0.577226, 0.5916324, 0.576326, 0.5790992, 
    0.5745099, 0.5704064, 0.5652554, 0.5557796, 0.5579705, 0.5500701, 
    0.6320087, 0.6270216, 0.6274614, 0.6222515, 0.6184042, 0.6100848, 
    0.5967935, 0.6017841, 0.5926306, 0.5907965, 0.6047065, 0.5961561, 
    0.6236895, 0.6192213, 0.6218816, 0.6316144, 0.6006317, 0.6164886, 
    0.5872829, 0.5958179, 0.5709909, 0.5833054, 0.5591773, 0.5489372, 
    0.539349, 0.5281939, 0.6243045, 0.6276891, 0.6216328, 0.6132728, 
    0.6055417, 0.5952963, 0.5942509, 0.5923365, 0.5873856, 0.58323, 
    0.5917304, 0.5821894, 0.6181839, 0.5992603, 0.6289686, 0.619988, 
    0.6137654, 0.6164945, 0.6023554, 0.5990334, 0.5855774, 0.5925251, 
    0.5514591, 0.5695391, 0.5197455, 0.5335408, 0.6288722, 0.6243168, 
    0.6085171, 0.6160236, 0.5946144, 0.5893707, 0.5851169, 0.5796882, 
    0.5791036, 0.5758937, 0.5811558, 0.5761018, 0.5952745, 0.5866885, 
    0.6103198, 0.6045479, 0.6072021, 0.6101155, 0.6011335, 0.591596, 
    0.5913944, 0.5883436, 0.5797637, 0.594528, 0.549133, 0.5770618, 
    0.6193573, 0.610616, 0.6093718, 0.6127528, 0.5898958, 0.5981546, 
    0.5759721, 0.5819481, 0.5721648, 0.5770212, 0.5777364, 0.5839904, 
    0.5878916, 0.597775, 0.6058449, 0.6122624, 0.610769, 0.6037242, 
    0.5910142, 0.5790499, 0.5816655, 0.572907, 0.5961608, 0.5863825, 
    0.5901568, 0.5803279, 0.6019165, 0.5835155, 0.6066403, 0.6046049, 
    0.5983188, 0.5857195, 0.5829432, 0.5799791, 0.581808, 0.5906927, 
    0.5921521, 0.5984718, 0.6002185, 0.6050481, 0.6090522, 0.6053931, 
    0.6015553, 0.5906897, 0.5809364, 0.5703478, 0.5677645, 0.5554627, 
    0.5654694, 0.5489781, 0.5629873, 0.5387954, 0.5824559, 0.5634043, 
    0.5980337, 0.5942801, 0.5875028, 0.5720325, 0.580374, 0.5706224, 
    0.5922094, 0.6034806, 0.6064069, 0.6118715, 0.6062822, 0.6067364, 
    0.6013978, 0.6031123, 0.5903297, 0.5971882, 0.5777539, 0.5706997, 
    0.5508961, 0.5388426, 0.5266474, 0.5212861, 0.5196574, 0.5189768,
  0.1245598, 0.1212654, 0.1219025, 0.1192703, 0.1207271, 0.1190085, 
    0.1238886, 0.1211354, 0.1228895, 0.1242617, 0.1142441, 0.1191536, 
    0.109257, 0.1123063, 0.1047288, 0.1097285, 0.1037353, 0.1048717, 
    0.1014719, 0.1024399, 0.0981542, 0.1010267, 0.09597109, 0.09883647, 
    0.09838513, 0.1011221, 0.1181577, 0.1148495, 0.1183551, 0.11788, 
    0.1180932, 0.1206968, 0.1220193, 0.1248138, 0.1243042, 0.122253, 
    0.1176668, 0.119214, 0.1153349, 0.1154218, 0.1111777, 0.1130813, 
    0.1060697, 0.1080391, 0.1023994, 0.1038029, 0.1024651, 0.1028698, 
    0.1024598, 0.1045223, 0.103636, 0.1054605, 0.1127234, 0.110563, 0.117069, 
    0.1210708, 0.1237671, 0.125698, 0.1254242, 0.1249028, 0.1222411, 
    0.1197649, 0.1178949, 0.1166522, 0.1154343, 0.1117862, 0.1098804, 
    0.1056735, 0.1064268, 0.1051525, 0.1039431, 0.1019285, 0.1022587, 
    0.1013761, 0.1051863, 0.1026457, 0.106857, 0.1056964, 0.1151028, 
    0.1187957, 0.1203818, 0.1217799, 0.1252138, 0.1228372, 0.1237713, 
    0.1215551, 0.1201571, 0.1208476, 0.1166183, 0.1182535, 0.109768, 
    0.1133836, 0.1040838, 0.106272, 0.1035629, 0.1049408, 0.1025855, 
    0.104704, 0.1010487, 0.1002616, 0.1007991, 0.09874305, 0.1048221, 
    0.1024649, 0.1208669, 0.1207541, 0.1202296, 0.1225437, 0.1226861, 
    0.1248277, 0.1229213, 0.1221138, 0.1200764, 0.1188792, 0.1177467, 
    0.115276, 0.1125478, 0.1087891, 0.1061294, 0.1043655, 0.1054454, 
    0.1044917, 0.1055581, 0.1060598, 0.1005561, 0.1036276, 0.09903741, 
    0.09928861, 0.1013551, 0.09926029, 0.120675, 0.1213244, 0.1235921, 
    0.1218157, 0.125062, 0.1232394, 0.1221974, 0.1182189, 0.117354, 
    0.1165544, 0.1149836, 0.1129834, 0.1095177, 0.1065475, 0.1038731, 
    0.1040678, 0.1039992, 0.1034061, 0.1048784, 0.1031654, 0.1028792, 
    0.1036282, 0.09932227, 0.1005427, 0.09929395, 0.1000876, 0.1211132, 
    0.1200225, 0.1206112, 0.1195053, 0.1202838, 0.1168412, 0.1158188, 
    0.111096, 0.1130226, 0.1099648, 0.1127101, 0.1122211, 0.1098652, 
    0.112561, 0.1067099, 0.1106587, 0.103383, 0.1072624, 0.1031424, 
    0.1038845, 0.1026574, 0.1015647, 0.1001989, 0.09770387, 0.09827874, 
    0.0962114, 0.1184059, 0.117008, 0.117131, 0.1156766, 0.1146068, 
    0.1123057, 0.1086645, 0.1100267, 0.107533, 0.1070358, 0.1108271, 
    0.108491, 0.1160774, 0.1148338, 0.1155736, 0.1182951, 0.1097116, 
    0.1140755, 0.1060857, 0.108399, 0.1017201, 0.1050138, 0.0985959, 
    0.09591629, 0.09343121, 0.09056965, 0.116249, 0.1171947, 0.1155043, 
    0.1131856, 0.1110563, 0.1082571, 0.1079729, 0.1074532, 0.1061134, 
    0.1049935, 0.1072889, 0.1047137, 0.1145457, 0.1093371, 0.117553, 
    0.1150468, 0.1133217, 0.1140771, 0.110183, 0.1092751, 0.1056256, 
    0.1075044, 0.09657379, 0.1013343, 0.08842358, 0.09193733, 0.117526, 
    0.1162524, 0.111874, 0.1139466, 0.1080717, 0.1066499, 0.1055015, 
    0.1040424, 0.1038857, 0.1030269, 0.1044361, 0.1030825, 0.1082512, 
    0.1059253, 0.1123705, 0.1107836, 0.1115123, 0.1123142, 0.1098487, 
    0.1072525, 0.1071978, 0.1063722, 0.1040628, 0.1080482, 0.09596737, 
    0.1033393, 0.1148715, 0.1124522, 0.1121093, 0.1130418, 0.106792, 
    0.1090354, 0.1030478, 0.1046489, 0.1020324, 0.1033283, 0.1035196, 
    0.1051981, 0.1062501, 0.1089319, 0.1111395, 0.1129064, 0.1124943, 
    0.1105579, 0.1070948, 0.1038713, 0.104573, 0.1022301, 0.1084923, 
    0.1058427, 0.1068626, 0.104214, 0.1100629, 0.1050704, 0.1113579, 
    0.1107993, 0.1090802, 0.1056639, 0.1049164, 0.1041204, 0.1046113, 
    0.1070077, 0.1074032, 0.1091219, 0.1095987, 0.1109208, 0.1120213, 
    0.1110155, 0.1099641, 0.1070069, 0.1043773, 0.1015491, 0.1008633, 
    0.09762087, 0.1002556, 0.09592704, 0.09959982, 0.09328857, 0.1047854, 
    0.0997098, 0.1090024, 0.1079808, 0.1061451, 0.1019972, 0.1042263, 
    0.1016221, 0.1074188, 0.1104911, 0.1112938, 0.1127985, 0.1112596, 
    0.1113843, 0.109921, 0.1103902, 0.1069094, 0.108772, 0.1035243, 
    0.1016427, 0.09642681, 0.09330068, 0.09017538, 0.08881354, 0.08840127, 
    0.08822922,
  0.008816513, 0.008483844, 0.008547862, 0.008284352, 0.008429865, 
    0.008258285, 0.008748401, 0.008470795, 0.008647338, 0.008786242, 
    0.007788455, 0.008272728, 0.007306031, 0.007599852, 0.006876457, 
    0.007351221, 0.006783308, 0.006889892, 0.006572567, 0.006662445, 
    0.006267461, 0.006531364, 0.006069169, 0.006329834, 0.00628855, 
    0.00654019, 0.008173742, 0.007847675, 0.00819333, 0.008146219, 
    0.008167345, 0.008426828, 0.008559614, 0.008842318, 0.008790549, 
    0.008583145, 0.008125095, 0.00827874, 0.007895251, 0.007903779, 
    0.007490678, 0.0076751, 0.007002808, 0.007189693, 0.006658677, 
    0.006789634, 0.006664784, 0.006702481, 0.006664294, 0.006857059, 
    0.006774012, 0.006945321, 0.007640325, 0.007431428, 0.008065974, 
    0.008464317, 0.008736094, 0.008932381, 0.008904455, 0.008851374, 
    0.008581941, 0.008333667, 0.00814769, 0.008024835, 0.007905005, 
    0.007549481, 0.007365801, 0.006965403, 0.007036582, 0.00691631, 
    0.006802758, 0.006614916, 0.006645594, 0.006563698, 0.006919489, 
    0.006681604, 0.007077337, 0.006967568, 0.0078725, 0.008237107, 
    0.008395303, 0.008535527, 0.008883022, 0.00864206, 0.008736522, 
    0.008512935, 0.008372835, 0.008441939, 0.008021493, 0.008183249, 
    0.00735501, 0.007704526, 0.006815937, 0.007021935, 0.00676718, 
    0.006896388, 0.006675994, 0.006874129, 0.006533403, 0.006460744, 
    0.006510335, 0.00632128, 0.006885224, 0.006664773, 0.008443874, 
    0.008432576, 0.008380086, 0.008612443, 0.008626803, 0.008843733, 
    0.008650547, 0.008569125, 0.008364772, 0.00824541, 0.008133008, 
    0.007889473, 0.007623275, 0.007261262, 0.007008455, 0.006842351, 
    0.006943893, 0.006854192, 0.006954514, 0.00700188, 0.006487897, 
    0.006773233, 0.006348239, 0.006371274, 0.006561754, 0.006368676, 
    0.00842465, 0.008489762, 0.00871837, 0.008539122, 0.008867574, 
    0.008682692, 0.008577542, 0.008179816, 0.008094142, 0.008015191, 
    0.007860808, 0.007665587, 0.007331005, 0.007048009, 0.006796196, 
    0.006814439, 0.006808012, 0.006752523, 0.006890517, 0.006730049, 
    0.006703356, 0.006773282, 0.006374363, 0.006486661, 0.006371764, 
    0.006444714, 0.008468565, 0.008359384, 0.008418261, 0.008307764, 
    0.008385498, 0.008043485, 0.007942784, 0.007482796, 0.007669391, 
    0.007373905, 0.00763903, 0.007591586, 0.007364342, 0.007624551, 
    0.007063393, 0.007440643, 0.006750372, 0.007115807, 0.006727901, 
    0.006797272, 0.006682689, 0.00658117, 0.006454966, 0.006226392, 
    0.006278829, 0.006090898, 0.008198375, 0.008059956, 0.008072106, 
    0.007928802, 0.007823912, 0.007599794, 0.007249357, 0.007379843, 
    0.007141515, 0.007094294, 0.007456861, 0.007232789, 0.007968214, 
    0.007846131, 0.007918687, 0.008187383, 0.007349601, 0.007771988, 
    0.007004323, 0.007224003, 0.006595577, 0.006903258, 0.006307818, 
    0.00606422, 0.005840987, 0.005587189, 0.007985102, 0.008078399, 
    0.007911881, 0.007685247, 0.00747896, 0.007210468, 0.007183382, 
    0.007133932, 0.007006941, 0.006901342, 0.007118321, 0.006875042, 
    0.007817945, 0.007313693, 0.008113837, 0.007867006, 0.007698496, 
    0.007772142, 0.007394862, 0.007307758, 0.006960886, 0.007138795, 
    0.006123717, 0.006559829, 0.005399156, 0.005708055, 0.008111161, 
    0.007985434, 0.007557976, 0.007759404, 0.007192792, 0.007057707, 
    0.00694918, 0.006812058, 0.006797382, 0.006717126, 0.006848974, 
    0.006722311, 0.007209904, 0.006989166, 0.007606071, 0.007452673, 
    0.00752299, 0.007600612, 0.007362757, 0.007114864, 0.007109669, 
    0.007031419, 0.006813976, 0.007190556, 0.006068842, 0.00674629, 
    0.007849822, 0.007614, 0.007580758, 0.007671264, 0.00707117, 0.007284815, 
    0.00671908, 0.006868951, 0.006624565, 0.006745254, 0.006763133, 
    0.006920598, 0.007019862, 0.007274918, 0.007486992, 0.007658098, 
    0.007618084, 0.007430928, 0.007099895, 0.006796036, 0.006861827, 
    0.006642929, 0.007232909, 0.006981374, 0.00707787, 0.006828134, 
    0.007383323, 0.00690859, 0.007508076, 0.007454178, 0.0072891, 
    0.006964504, 0.006894088, 0.006819366, 0.006865417, 0.00709163, 
    0.007129181, 0.007293092, 0.00733877, 0.007465893, 0.00757223, 
    0.007475025, 0.007373836, 0.00709155, 0.006843453, 0.006579727, 
    0.006516266, 0.006218839, 0.006460192, 0.006065197, 0.006399859, 
    0.00582826, 0.006881786, 0.006409961, 0.00728166, 0.007184137, 
    0.007009942, 0.006621301, 0.006829295, 0.006586495, 0.007130658, 
    0.007424506, 0.007501886, 0.007647614, 0.007498577, 0.007510627, 
    0.007369694, 0.00741479, 0.007082305, 0.007259628, 0.006763572, 
    0.006588399, 0.006110398, 0.005829336, 0.005552492, 0.005433173, 
    0.005397211, 0.005382224,
  0.0001783862, 0.000169057, 0.0001708417, 0.0001635287, 0.0001675562, 
    0.00016281, 0.000176465, 0.0001686939, 0.0001736249, 0.0001775317, 
    0.0001500069, 0.0001632081, 0.0001371637, 0.0001449485, 0.0001259969, 
    0.0001383534, 0.0001236099, 0.0001263422, 0.0001182561, 0.0001205315, 
    0.0001106214, 0.0001172169, 0.0001057351, 0.0001121708, 0.0001111446, 
    0.0001174393, 0.0001604851, 0.0001516049, 0.000161023, 0.0001597302, 
    0.0001603096, 0.0001674719, 0.0001711699, 0.0001791155, 0.0001776532, 
    0.0001718275, 0.0001591515, 0.0001633738, 0.0001528918, 0.0001531228, 
    0.0001420423, 0.0001469609, 0.0001292544, 0.000134114, 0.0001204358, 
    0.0001237716, 0.0001205908, 0.0001215488, 0.0001205784, 0.0001254987, 
    0.0001233724, 0.0001277695, 0.0001460299, 0.0001404717, 0.0001575348, 
    0.0001685138, 0.0001761185, 0.0001816673, 0.0001808751, 0.0001793717, 
    0.0001717938, 0.0001648906, 0.0001597705, 0.0001564125, 0.000153156, 
    0.0001436057, 0.0001387378, 0.0001282877, 0.000130129, 0.0001270219, 
    0.0001241073, 0.0001193267, 0.000120104, 0.0001180322, 0.0001271037, 
    0.0001210181, 0.0001311865, 0.0001283436, 0.0001522761, 0.0001622267, 
    0.0001665972, 0.0001704974, 0.0001802676, 0.0001734769, 0.0001761305, 
    0.0001698673, 0.0001659745, 0.0001678916, 0.0001563215, 0.0001607461, 
    0.0001384533, 0.00014775, 0.0001244446, 0.0001297495, 0.0001231979, 
    0.0001265092, 0.0001208755, 0.000125937, 0.0001172683, 0.0001154418, 
    0.0001166876, 0.0001119579, 0.0001262221, 0.0001205906, 0.0001679453, 
    0.0001676315, 0.0001661753, 0.0001726472, 0.0001730493, 0.0001791555, 
    0.0001737148, 0.0001714355, 0.0001657512, 0.0001624553, 0.0001593682, 
    0.0001527353, 0.0001455741, 0.0001359879, 0.0001294005, 0.0001251214, 
    0.0001277326, 0.0001254252, 0.0001280066, 0.0001292304, 0.0001161234, 
    0.0001233525, 0.0001126291, 0.0001132034, 0.0001179831, 0.0001131386, 
    0.0001674114, 0.0001692217, 0.0001756197, 0.0001705977, 0.0001798301, 
    0.000174617, 0.0001716708, 0.0001606519, 0.0001583045, 0.0001561498, 
    0.0001519597, 0.0001467061, 0.0001378208, 0.0001304253, 0.0001239394, 
    0.0001244062, 0.0001242417, 0.0001228238, 0.0001263582, 0.0001222508, 
    0.0001215711, 0.0001233537, 0.0001132805, 0.0001160924, 0.0001132156, 
    0.0001150398, 0.0001686318, 0.000165602, 0.000167234, 0.0001641748, 
    0.0001663254, 0.0001569211, 0.0001541808, 0.0001418331, 0.000146808, 
    0.0001389516, 0.0001459953, 0.0001447279, 0.0001386994, 0.0001456082, 
    0.0001308245, 0.0001407158, 0.0001227689, 0.000132187, 0.000122196, 
    0.0001239669, 0.0001210456, 0.0001184734, 0.0001152968, 0.0001096044, 
    0.0001109033, 0.0001062675, 0.0001611615, 0.0001573705, 0.0001577023, 
    0.0001538012, 0.0001509629, 0.0001449469, 0.0001356757, 0.0001391083, 
    0.0001328565, 0.0001316272, 0.0001411453, 0.0001352416, 0.0001548715, 
    0.000151563, 0.0001535269, 0.0001608596, 0.0001383107, 0.0001495632, 
    0.0001292936, 0.0001350114, 0.0001188375, 0.0001266859, 0.0001116232, 
    0.0001056139, 0.0001001878, 9.411546e-05, 0.0001553307, 0.0001578742, 
    0.0001533424, 0.0001472329, 0.0001417313, 0.0001346572, 0.0001339491, 
    0.0001326589, 0.0001293613, 0.0001266366, 0.0001322524, 0.0001259605, 
    0.0001508021, 0.0001373652, 0.0001588433, 0.0001521274, 0.0001475882, 
    0.0001495673, 0.0001395049, 0.0001372091, 0.0001281711, 0.0001327856, 
    0.0001070732, 0.0001179346, 8.968443e-05, 9.699433e-05, 0.00015877, 
    0.0001553397, 0.0001438319, 0.0001492245, 0.000134195, 0.0001306769, 
    0.000127869, 0.0001243453, 0.0001239697, 0.0001219216, 0.0001252913, 
    0.0001220536, 0.0001346425, 0.0001289016, 0.0001451145, 0.0001410343, 
    0.0001429007, 0.0001449688, 0.0001386575, 0.0001321624, 0.0001320271, 
    0.0001299952, 0.0001243945, 0.0001341365, 0.0001057272, 0.0001226649, 
    0.0001516627, 0.0001453263, 0.000144439, 0.0001468581, 0.0001310264, 
    0.0001366061, 0.0001219713, 0.000125804, 0.000119571, 0.0001226384, 
    0.0001230945, 0.0001271323, 0.0001296958, 0.0001363463, 0.0001419444, 
    0.0001465055, 0.0001454354, 0.0001404585, 0.0001317729, 0.0001239353, 
    0.0001256211, 0.0001200364, 0.0001352447, 0.0001287002, 0.0001312004, 
    0.000124757, 0.0001392002, 0.0001268233, 0.0001425043, 0.0001410742, 
    0.0001367187, 0.0001282645, 0.00012645, 0.0001245324, 0.0001257133, 
    0.000131558, 0.0001325351, 0.0001368236, 0.0001380253, 0.0001413847, 
    0.0001442117, 0.0001416268, 0.0001389498, 0.0001315559, 0.0001251497, 
    0.0001184369, 0.0001168368, 0.0001094177, 0.000115428, 0.0001056379, 
    0.0001139174, 9.988096e-05, 0.0001261338, 0.0001141699, 0.0001365233, 
    0.0001339688, 0.0001294391, 0.0001194884, 0.0001247868, 0.000118608, 
    0.0001325736, 0.0001402886, 0.0001423398, 0.0001462249, 0.000142252, 
    0.0001425721, 0.0001388404, 0.0001400316, 0.0001313156, 0.000135945, 
    0.0001231058, 0.0001186561, 0.000106746, 9.990684e-05, 9.329336e-05, 
    9.048166e-05, 8.963887e-05, 8.92883e-05,
  1.137658e-06, 1.055336e-06, 1.070966e-06, 1.007284e-06, 1.042236e-06, 
    1.001078e-06, 1.120581e-06, 1.052163e-06, 1.095453e-06, 1.130054e-06, 
    8.921508e-07, 1.004515e-06, 7.861224e-07, 8.4999e-07, 6.967555e-07, 
    7.958017e-07, 6.780116e-07, 6.994771e-07, 6.364473e-07, 6.540302e-07, 
    5.783602e-07, 6.284581e-07, 5.419437e-07, 5.900326e-07, 5.82295e-07, 
    6.301658e-07, 9.810678e-07, 9.055746e-07, 9.856882e-07, 9.745924e-07, 
    9.795609e-07, 1.041502e-06, 1.073847e-06, 1.144157e-06, 1.131135e-06, 
    1.079623e-06, 9.69635e-07, 1.005946e-06, 9.164206e-07, 9.183711e-07, 
    8.260006e-07, 8.667017e-07, 7.225425e-07, 7.614464e-07, 6.532889e-07, 
    6.792768e-07, 6.544908e-07, 6.619313e-07, 6.543943e-07, 6.928328e-07, 
    6.76153e-07, 7.107579e-07, 8.589606e-07, 8.131089e-07, 9.558203e-07, 
    1.05059e-06, 1.117508e-06, 1.166969e-06, 1.159875e-06, 1.146442e-06, 
    1.079327e-06, 1.01907e-06, 9.749374e-07, 9.462589e-07, 9.186518e-07, 
    8.388851e-07, 7.989353e-07, 7.148651e-07, 7.295059e-07, 7.048439e-07, 
    6.81906e-07, 6.447057e-07, 6.507175e-07, 6.34724e-07, 7.054904e-07, 
    6.578064e-07, 7.379483e-07, 7.15308e-07, 9.112282e-07, 9.960484e-07, 
    1.033888e-06, 1.067946e-06, 1.154443e-06, 1.094148e-06, 1.117615e-06, 
    1.062425e-06, 1.028475e-06, 1.04516e-06, 9.454841e-07, 9.83309e-07, 
    7.966151e-07, 8.732765e-07, 6.845509e-07, 7.264824e-07, 6.747887e-07, 
    7.007947e-07, 6.566997e-07, 6.962835e-07, 6.288527e-07, 6.148704e-07, 
    6.243983e-07, 5.884252e-07, 6.985306e-07, 6.544888e-07, 1.045629e-06, 
    1.042892e-06, 1.03022e-06, 1.086836e-06, 1.090378e-06, 1.144514e-06, 
    1.096247e-06, 1.076179e-06, 1.026535e-06, 9.980189e-07, 9.714904e-07, 
    9.151002e-07, 8.551771e-07, 7.765853e-07, 7.237046e-07, 6.898653e-07, 
    7.104661e-07, 6.922538e-07, 7.126366e-07, 7.223513e-07, 6.200792e-07, 
    6.759977e-07, 5.934967e-07, 5.978453e-07, 6.343466e-07, 5.973541e-07, 
    1.040974e-06, 1.056776e-06, 1.113088e-06, 1.068825e-06, 1.150534e-06, 
    1.104215e-06, 1.078247e-06, 9.825001e-07, 9.623909e-07, 9.44024e-07, 
    9.08561e-07, 8.64581e-07, 7.914643e-07, 7.31869e-07, 6.805907e-07, 
    6.842499e-07, 6.829597e-07, 6.718664e-07, 6.996036e-07, 6.673965e-07, 
    6.621048e-07, 6.760072e-07, 5.984294e-07, 6.198414e-07, 5.97938e-07, 
    6.118041e-07, 1.05162e-06, 1.02524e-06, 1.039429e-06, 1.012872e-06, 
    1.031523e-06, 9.505888e-07, 9.273175e-07, 8.242809e-07, 8.654288e-07, 
    8.006792e-07, 8.586729e-07, 8.481631e-07, 7.986221e-07, 8.554592e-07, 
    7.350558e-07, 8.151089e-07, 6.714381e-07, 7.459585e-07, 6.669699e-07, 
    6.808062e-07, 6.580202e-07, 6.381213e-07, 6.13764e-07, 5.707305e-07, 
    5.804793e-07, 5.458821e-07, 9.868794e-07, 9.544192e-07, 9.572485e-07, 
    9.241054e-07, 9.001752e-07, 8.499769e-07, 7.740578e-07, 8.019578e-07, 
    7.513304e-07, 7.414739e-07, 8.186312e-07, 7.705468e-07, 9.331696e-07, 
    9.052219e-07, 9.217857e-07, 9.842846e-07, 7.954533e-07, 8.884324e-07, 
    7.228541e-07, 7.686874e-07, 6.409287e-07, 7.021903e-07, 5.859002e-07, 
    5.410488e-07, 5.013538e-07, 4.578789e-07, 9.37065e-07, 9.58716e-07, 
    9.20226e-07, 8.68967e-07, 8.234437e-07, 7.658275e-07, 7.601179e-07, 
    7.497439e-07, 7.233927e-07, 7.018006e-07, 7.464825e-07, 6.964682e-07, 
    8.988242e-07, 7.877594e-07, 9.669975e-07, 9.099742e-07, 8.719275e-07, 
    8.884664e-07, 8.051972e-07, 7.864904e-07, 7.139404e-07, 7.50761e-07, 
    5.518563e-07, 6.339734e-07, 4.268141e-07, 4.783626e-07, 9.663707e-07, 
    9.371415e-07, 8.407526e-07, 8.85596e-07, 7.620992e-07, 7.338766e-07, 
    7.115461e-07, 6.837722e-07, 6.808284e-07, 6.648323e-07, 6.912007e-07, 
    6.658603e-07, 7.657083e-07, 7.197379e-07, 8.513654e-07, 8.177208e-07, 
    8.330686e-07, 8.501578e-07, 7.982794e-07, 7.457611e-07, 7.446768e-07, 
    7.284398e-07, 6.841593e-07, 7.616281e-07, 5.418861e-07, 6.706275e-07, 
    9.060604e-07, 8.531218e-07, 8.457723e-07, 8.658462e-07, 7.366684e-07, 
    7.815957e-07, 6.652195e-07, 6.952359e-07, 6.465938e-07, 6.704191e-07, 
    6.739813e-07, 7.057162e-07, 7.260549e-07, 7.794885e-07, 8.251957e-07, 
    8.629129e-07, 8.540255e-07, 8.130004e-07, 7.426405e-07, 6.80559e-07, 
    6.937961e-07, 6.501942e-07, 7.705717e-07, 7.181387e-07, 7.380595e-07, 
    6.870027e-07, 8.02708e-07, 7.032755e-07, 8.298026e-07, 8.180477e-07, 
    7.825088e-07, 7.146814e-07, 7.003281e-07, 6.852399e-07, 6.945212e-07, 
    7.409199e-07, 7.487506e-07, 7.833598e-07, 7.931286e-07, 8.205964e-07, 
    8.438914e-07, 8.225855e-07, 8.006643e-07, 7.409029e-07, 6.900877e-07, 
    6.378405e-07, 6.25542e-07, 5.693333e-07, 6.147654e-07, 5.412268e-07, 
    6.032639e-07, 4.99133e-07, 6.97835e-07, 6.051819e-07, 7.809235e-07, 
    7.602767e-07, 7.240114e-07, 6.459557e-07, 6.872363e-07, 6.391589e-07, 
    7.490592e-07, 8.11609e-07, 8.284489e-07, 8.605805e-07, 8.277256e-07, 
    8.303608e-07, 7.997718e-07, 8.095043e-07, 7.389806e-07, 7.762376e-07, 
    6.740692e-07, 6.395296e-07, 5.49428e-07, 4.9932e-07, 4.520723e-07, 
    4.32361e-07, 4.264976e-07, 4.240648e-07,
  1.368999e-09, 1.195315e-09, 1.227759e-09, 1.097192e-09, 1.16832e-09, 
    1.084703e-09, 1.332409e-09, 1.18876e-09, 1.279097e-09, 1.352671e-09, 
    8.726678e-10, 1.091613e-09, 6.804365e-10, 7.944576e-10, 5.306708e-10, 
    6.973585e-10, 5.008224e-10, 5.350512e-10, 4.367149e-10, 4.634763e-10, 
    3.522443e-10, 4.247332e-10, 3.025752e-10, 3.68715e-10, 3.577673e-10, 
    4.272849e-10, 1.044722e-09, 8.980371e-10, 1.053913e-09, 1.03188e-09, 
    1.041729e-09, 1.166811e-09, 1.233768e-09, 1.382997e-09, 1.354987e-09, 
    1.24584e-09, 1.022082e-09, 1.094495e-09, 9.186933e-10, 9.224236e-10, 
    7.509838e-10, 8.251866e-10, 5.726469e-10, 6.37898e-10, 4.623373e-10, 
    5.028187e-10, 4.641846e-10, 4.756741e-10, 4.640361e-10, 5.243768e-10, 
    4.978936e-10, 5.533347e-10, 8.109078e-10, 7.27939e-10, 9.949231e-10, 
    1.185516e-09, 1.325855e-09, 1.43246e-09, 1.417024e-09, 1.38793e-09, 
    1.24522e-09, 1.121028e-09, 1.032563e-09, 9.762555e-10, 9.229608e-10, 
    7.742399e-10, 7.028647e-10, 5.600413e-10, 5.841588e-10, 5.437247e-10, 
    5.069766e-10, 4.492179e-10, 4.583937e-10, 4.341212e-10, 5.447722e-10, 
    4.692932e-10, 5.982146e-10, 5.607657e-10, 9.087879e-10, 1.074611e-09, 
    1.151212e-09, 1.221471e-09, 1.405237e-09, 1.276345e-09, 1.326083e-09, 
    1.209999e-09, 1.140157e-09, 1.174328e-09, 9.747475e-10, 1.049177e-09, 
    6.987861e-10, 8.373749e-10, 5.111707e-10, 5.791513e-10, 4.957474e-10, 
    5.371762e-10, 4.675858e-10, 5.299115e-10, 4.253224e-10, 4.046165e-10, 
    4.186881e-10, 3.664311e-10, 5.335261e-10, 4.641816e-10, 1.175293e-09, 
    1.169667e-09, 1.143717e-09, 1.260961e-09, 1.268407e-09, 1.383768e-09, 
    1.280771e-09, 1.238638e-09, 1.136205e-09, 1.078561e-09, 1.025745e-09, 
    9.161709e-10, 8.039571e-10, 6.638923e-10, 5.745629e-10, 5.19632e-10, 
    5.528589e-10, 5.234497e-10, 5.563988e-10, 5.723316e-10, 4.122892e-10, 
    4.976492e-10, 3.73653e-10, 3.798838e-10, 4.335539e-10, 3.791782e-10, 
    1.165729e-09, 1.198293e-09, 1.316445e-09, 1.223301e-09, 1.396775e-09, 
    1.297615e-09, 1.24296e-09, 1.047569e-09, 1.007812e-09, 9.719078e-10, 
    9.037087e-10, 8.212672e-10, 6.897589e-10, 5.880826e-10, 5.048951e-10, 
    5.106926e-10, 5.08646e-10, 4.911609e-10, 5.35255e-10, 4.841729e-10, 
    4.759433e-10, 4.976639e-10, 3.807236e-10, 4.119375e-10, 3.80017e-10, 
    4.001224e-10, 1.187638e-09, 1.133568e-09, 1.162559e-09, 1.108474e-09, 
    1.146379e-09, 9.846967e-10, 9.395932e-10, 7.478974e-10, 8.228337e-10, 
    7.059344e-10, 8.103785e-10, 7.911202e-10, 7.023142e-10, 8.044742e-10, 
    5.933876e-10, 7.315001e-10, 4.904899e-10, 6.116515e-10, 4.835077e-10, 
    5.052359e-10, 4.696228e-10, 4.392398e-10, 4.029928e-10, 3.416196e-10, 
    3.552145e-10, 3.078175e-10, 1.056287e-09, 9.921811e-10, 9.977202e-10, 
    9.33417e-10, 8.878042e-10, 7.944333e-10, 6.595292e-10, 7.081877e-10, 
    6.207141e-10, 6.041166e-10, 7.377826e-10, 6.534844e-10, 9.508747e-10, 
    8.973662e-10, 9.289654e-10, 1.051119e-09, 6.967466e-10, 8.656784e-10, 
    5.731605e-10, 6.502898e-10, 4.43485e-10, 5.394307e-10, 3.628538e-10, 
    3.013888e-10, 2.504595e-10, 1.987538e-10, 9.584068e-10, 1.000597e-09, 
    9.259754e-10, 8.293805e-10, 7.463953e-10, 6.453865e-10, 6.356327e-10, 
    6.18033e-10, 5.740483e-10, 5.388004e-10, 6.125331e-10, 5.302084e-10, 
    8.852516e-10, 6.832888e-10, 1.016879e-09, 9.063987e-10, 8.348698e-10, 
    8.657418e-10, 7.139077e-10, 6.810766e-10, 5.585289e-10, 6.197514e-10, 
    3.158315e-10, 4.329933e-10, 1.646376e-10, 2.225616e-10, 1.015644e-09, 
    9.585547e-10, 7.776276e-10, 8.603589e-10, 6.39012e-10, 5.914224e-10, 
    5.546192e-10, 5.099348e-10, 5.05271e-10, 4.801792e-10, 5.217654e-10, 
    4.817788e-10, 6.451824e-10, 5.680313e-10, 7.969726e-10, 7.361571e-10, 
    7.637128e-10, 7.94764e-10, 7.0171e-10, 6.113186e-10, 6.09494e-10, 
    5.823917e-10, 5.10551e-10, 6.382079e-10, 3.025e-10, 4.892226e-10, 
    8.98957e-10, 8.001894e-10, 7.86759e-10, 8.236047e-10, 5.96077e-10, 
    6.725674e-10, 4.807816e-10, 5.282292e-10, 4.520929e-10, 4.888946e-10, 
    4.944788e-10, 5.451383e-10, 5.784443e-10, 6.689146e-10, 7.495386e-10, 
    8.181881e-10, 8.018445e-10, 7.27746e-10, 6.060737e-10, 5.048453e-10, 
    5.259203e-10, 4.575924e-10, 6.535268e-10, 5.654051e-10, 5.984011e-10, 
    5.150688e-10, 7.095113e-10, 5.411868e-10, 7.578225e-10, 7.367405e-10, 
    6.741522e-10, 5.59741e-10, 5.364232e-10, 5.122653e-10, 5.270825e-10, 
    6.031883e-10, 6.16356e-10, 6.756303e-10, 6.926714e-10, 7.412957e-10, 
    7.833333e-10, 7.448572e-10, 7.059081e-10, 6.031595e-10, 5.199874e-10, 
    4.38816e-10, 4.203881e-10, 3.396869e-10, 4.044629e-10, 3.016257e-10, 
    3.876996e-10, 2.477131e-10, 5.324075e-10, 3.904774e-10, 6.714011e-10, 
    6.359033e-10, 5.750696e-10, 4.511212e-10, 5.154405e-10, 4.408076e-10, 
    6.168769e-10, 7.252728e-10, 7.553855e-10, 8.138893e-10, 7.54084e-10, 
    7.588284e-10, 7.043359e-10, 7.215353e-10, 5.999409e-10, 6.632911e-10, 
    4.946169e-10, 4.41368e-10, 3.125651e-10, 2.479433e-10, 1.921904e-10, 
    1.705469e-10, 1.643027e-10, 1.617386e-10,
  4.068484e-13, 4.060851e-13, 4.062277e-13, 4.056534e-13, 4.059664e-13, 
    4.055985e-13, 4.066877e-13, 4.060563e-13, 4.064534e-13, 4.067767e-13, 
    4.046644e-13, 4.056289e-13, 4.038161e-13, 4.043195e-13, 4.031539e-13, 
    4.038908e-13, 4.030218e-13, 4.031733e-13, 4.027379e-13, 4.028564e-13, 
    4.023633e-13, 4.026848e-13, 4.021428e-13, 4.024364e-13, 4.023878e-13, 
    4.026961e-13, 4.054225e-13, 4.047763e-13, 4.054629e-13, 4.053659e-13, 
    4.054093e-13, 4.059597e-13, 4.062542e-13, 4.069099e-13, 4.067869e-13, 
    4.063072e-13, 4.053228e-13, 4.056416e-13, 4.048673e-13, 4.048838e-13, 
    4.041276e-13, 4.044551e-13, 4.033396e-13, 4.036281e-13, 4.028514e-13, 
    4.030306e-13, 4.028595e-13, 4.029105e-13, 4.028589e-13, 4.03126e-13, 
    4.030088e-13, 4.032542e-13, 4.043921e-13, 4.040259e-13, 4.052032e-13, 
    4.06042e-13, 4.066589e-13, 4.071271e-13, 4.070593e-13, 4.069316e-13, 
    4.063045e-13, 4.057583e-13, 4.053689e-13, 4.05121e-13, 4.048861e-13, 
    4.042303e-13, 4.039152e-13, 4.032839e-13, 4.033905e-13, 4.032117e-13, 
    4.03049e-13, 4.027933e-13, 4.028339e-13, 4.027264e-13, 4.032163e-13, 
    4.028822e-13, 4.034527e-13, 4.032871e-13, 4.048237e-13, 4.05554e-13, 
    4.058911e-13, 4.062001e-13, 4.070076e-13, 4.064413e-13, 4.066599e-13, 
    4.061497e-13, 4.058425e-13, 4.059928e-13, 4.051143e-13, 4.054421e-13, 
    4.038971e-13, 4.045088e-13, 4.030676e-13, 4.033684e-13, 4.029993e-13, 
    4.031827e-13, 4.028746e-13, 4.031505e-13, 4.026874e-13, 4.025956e-13, 
    4.02658e-13, 4.024262e-13, 4.031665e-13, 4.028595e-13, 4.05997e-13, 
    4.059723e-13, 4.058581e-13, 4.063737e-13, 4.064064e-13, 4.069133e-13, 
    4.064608e-13, 4.062756e-13, 4.058251e-13, 4.055714e-13, 4.053389e-13, 
    4.048562e-13, 4.043614e-13, 4.03743e-13, 4.033481e-13, 4.03105e-13, 
    4.032521e-13, 4.03122e-13, 4.032678e-13, 4.033382e-13, 4.026296e-13, 
    4.030077e-13, 4.024583e-13, 4.024859e-13, 4.027239e-13, 4.024828e-13, 
    4.05955e-13, 4.060982e-13, 4.066175e-13, 4.062081e-13, 4.069704e-13, 
    4.065348e-13, 4.062946e-13, 4.05435e-13, 4.052599e-13, 4.051018e-13, 
    4.048013e-13, 4.044378e-13, 4.038573e-13, 4.034079e-13, 4.030398e-13, 
    4.030655e-13, 4.030564e-13, 4.02979e-13, 4.031742e-13, 4.029481e-13, 
    4.029116e-13, 4.030078e-13, 4.024896e-13, 4.02628e-13, 4.024865e-13, 
    4.025757e-13, 4.060513e-13, 4.058135e-13, 4.05941e-13, 4.057031e-13, 
    4.058698e-13, 4.051581e-13, 4.049594e-13, 4.04114e-13, 4.044447e-13, 
    4.039287e-13, 4.043897e-13, 4.043048e-13, 4.039127e-13, 4.043637e-13, 
    4.034314e-13, 4.040416e-13, 4.02976e-13, 4.035121e-13, 4.029451e-13, 
    4.030413e-13, 4.028836e-13, 4.02749e-13, 4.025884e-13, 4.023162e-13, 
    4.023765e-13, 4.021661e-13, 4.054734e-13, 4.051911e-13, 4.052155e-13, 
    4.049322e-13, 4.047312e-13, 4.043194e-13, 4.037237e-13, 4.039387e-13, 
    4.035522e-13, 4.034788e-13, 4.040693e-13, 4.03697e-13, 4.050091e-13, 
    4.047733e-13, 4.049126e-13, 4.054506e-13, 4.038881e-13, 4.046336e-13, 
    4.033419e-13, 4.036829e-13, 4.027679e-13, 4.031927e-13, 4.024104e-13, 
    4.021376e-13, 4.019112e-13, 4.016812e-13, 4.050423e-13, 4.052282e-13, 
    4.048994e-13, 4.044735e-13, 4.041074e-13, 4.036612e-13, 4.036181e-13, 
    4.035403e-13, 4.033458e-13, 4.031899e-13, 4.03516e-13, 4.031519e-13, 
    4.047199e-13, 4.038287e-13, 4.052999e-13, 4.048131e-13, 4.044978e-13, 
    4.046339e-13, 4.039639e-13, 4.038189e-13, 4.032772e-13, 4.035479e-13, 
    4.022017e-13, 4.027214e-13, 4.015293e-13, 4.017871e-13, 4.052945e-13, 
    4.05043e-13, 4.042452e-13, 4.046102e-13, 4.03633e-13, 4.034227e-13, 
    4.032599e-13, 4.030621e-13, 4.030415e-13, 4.029304e-13, 4.031145e-13, 
    4.029375e-13, 4.036603e-13, 4.033192e-13, 4.043306e-13, 4.040622e-13, 
    4.041838e-13, 4.043208e-13, 4.039101e-13, 4.035106e-13, 4.035026e-13, 
    4.033827e-13, 4.030648e-13, 4.036295e-13, 4.021425e-13, 4.029704e-13, 
    4.047803e-13, 4.043448e-13, 4.042855e-13, 4.044481e-13, 4.034432e-13, 
    4.037813e-13, 4.029331e-13, 4.031431e-13, 4.02806e-13, 4.02969e-13, 
    4.029937e-13, 4.032179e-13, 4.033652e-13, 4.037652e-13, 4.041212e-13, 
    4.044242e-13, 4.043521e-13, 4.04025e-13, 4.034874e-13, 4.030396e-13, 
    4.031329e-13, 4.028304e-13, 4.036972e-13, 4.033076e-13, 4.034535e-13, 
    4.030848e-13, 4.039445e-13, 4.032004e-13, 4.041578e-13, 4.040647e-13, 
    4.037883e-13, 4.032825e-13, 4.031794e-13, 4.030724e-13, 4.03138e-13, 
    4.034747e-13, 4.035329e-13, 4.037949e-13, 4.038701e-13, 4.040849e-13, 
    4.042704e-13, 4.041006e-13, 4.039286e-13, 4.034746e-13, 4.031066e-13, 
    4.027472e-13, 4.026655e-13, 4.023076e-13, 4.025949e-13, 4.021386e-13, 
    4.025206e-13, 4.01899e-13, 4.031616e-13, 4.025329e-13, 4.037762e-13, 
    4.036193e-13, 4.033503e-13, 4.028017e-13, 4.030865e-13, 4.02756e-13, 
    4.035352e-13, 4.040141e-13, 4.04147e-13, 4.044052e-13, 4.041413e-13, 
    4.041622e-13, 4.039217e-13, 4.039976e-13, 4.034603e-13, 4.037403e-13, 
    4.029943e-13, 4.027585e-13, 4.021872e-13, 4.019e-13, 4.01652e-13, 
    4.015556e-13, 4.015278e-13, 4.015163e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 
    8.949648e-07, 8.94965e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 
    8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949647e-07, 
    8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.94965e-07, 8.949649e-07, 8.94965e-07, 8.949649e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 
    8.94965e-07, 8.949649e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 
    8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949649e-07, 
    8.94965e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 8.949649e-07, 
    8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949649e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 8.94965e-07, 
    8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.949646e-07, 8.949647e-07, 8.949647e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 
    8.949647e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.949649e-07, 8.949649e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.949646e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 
    8.949649e-07, 8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949649e-07, 
    8.949649e-07, 8.949649e-07, 8.94965e-07, 8.949648e-07, 8.949648e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 
    8.949646e-07, 8.949645e-07, 8.949644e-07, 8.949649e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949648e-07, 8.949648e-07, 8.949649e-07, 8.949649e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949646e-07, 8.949646e-07, 8.949644e-07, 8.949644e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949646e-07, 8.949647e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 
    8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.949645e-07, 8.949647e-07, 8.949646e-07, 8.949648e-07, 
    8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 
    8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949645e-07, 8.949644e-07, 
    8.949644e-07, 8.949644e-07, 8.949644e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.968902e-16, 6.986648e-16, 6.983201e-16, 6.9975e-16, 6.989572e-16, 
    6.998931e-16, 6.972505e-16, 6.987349e-16, 6.977876e-16, 6.970505e-16, 
    7.025202e-16, 6.998138e-16, 7.053292e-16, 7.036064e-16, 7.079312e-16, 
    7.050609e-16, 7.085094e-16, 7.078491e-16, 7.098371e-16, 7.092679e-16, 
    7.118062e-16, 7.100997e-16, 7.131213e-16, 7.113992e-16, 7.116685e-16, 
    7.100433e-16, 7.003595e-16, 7.021834e-16, 7.002512e-16, 7.005114e-16, 
    7.003948e-16, 6.989733e-16, 6.982561e-16, 6.967549e-16, 6.970277e-16, 
    6.981304e-16, 7.006285e-16, 6.997814e-16, 7.019166e-16, 7.018685e-16, 
    7.042418e-16, 7.031722e-16, 7.071561e-16, 7.06025e-16, 7.092916e-16, 
    7.084707e-16, 7.09253e-16, 7.090159e-16, 7.092561e-16, 7.080519e-16, 
    7.085679e-16, 7.075081e-16, 7.033724e-16, 7.045888e-16, 7.009576e-16, 
    6.987691e-16, 6.973155e-16, 6.962826e-16, 6.964286e-16, 6.967069e-16, 
    6.981369e-16, 6.994808e-16, 7.005039e-16, 7.011878e-16, 7.018616e-16, 
    7.038972e-16, 7.04975e-16, 7.073844e-16, 7.069504e-16, 7.076859e-16, 
    7.083891e-16, 7.09568e-16, 7.093741e-16, 7.098931e-16, 7.076669e-16, 
    7.091466e-16, 7.06703e-16, 7.073717e-16, 7.020425e-16, 7.000101e-16, 
    6.991435e-16, 6.983863e-16, 6.965409e-16, 6.978154e-16, 6.973131e-16, 
    6.985084e-16, 6.992671e-16, 6.98892e-16, 7.012065e-16, 7.00307e-16, 
    7.050389e-16, 7.030025e-16, 7.083071e-16, 7.070395e-16, 7.086108e-16, 
    7.078093e-16, 7.091821e-16, 7.079467e-16, 7.100865e-16, 7.105517e-16, 
    7.102337e-16, 7.114555e-16, 7.078781e-16, 7.092528e-16, 6.988814e-16, 
    6.989425e-16, 6.992278e-16, 6.979736e-16, 6.97897e-16, 6.967473e-16, 
    6.977705e-16, 6.982058e-16, 6.993112e-16, 6.999644e-16, 7.005851e-16, 
    7.01949e-16, 7.034705e-16, 7.055961e-16, 7.071217e-16, 7.081433e-16, 
    7.075171e-16, 7.0807e-16, 7.074518e-16, 7.071621e-16, 7.103773e-16, 
    7.085726e-16, 7.112799e-16, 7.111303e-16, 7.099054e-16, 7.111471e-16, 
    6.989855e-16, 6.986334e-16, 6.974096e-16, 6.983674e-16, 6.966221e-16, 
    6.97599e-16, 6.981603e-16, 7.003254e-16, 7.008012e-16, 7.012416e-16, 
    7.021115e-16, 7.032269e-16, 7.051816e-16, 7.068805e-16, 7.0843e-16, 
    7.083166e-16, 7.083565e-16, 7.087022e-16, 7.078454e-16, 7.088429e-16, 
    7.0901e-16, 7.085727e-16, 7.111102e-16, 7.103857e-16, 7.111271e-16, 
    7.106555e-16, 6.987479e-16, 6.993404e-16, 6.990202e-16, 6.996222e-16, 
    6.99198e-16, 7.010827e-16, 7.016473e-16, 7.042871e-16, 7.032048e-16, 
    7.049276e-16, 7.033801e-16, 7.036543e-16, 7.049828e-16, 7.034639e-16, 
    7.067864e-16, 7.045339e-16, 7.087156e-16, 7.064683e-16, 7.088563e-16, 
    7.084233e-16, 7.091404e-16, 7.097821e-16, 7.105893e-16, 7.12077e-16, 
    7.117328e-16, 7.129764e-16, 7.002236e-16, 7.009911e-16, 7.009239e-16, 
    7.017271e-16, 7.023208e-16, 7.036071e-16, 7.056675e-16, 7.048932e-16, 
    7.063149e-16, 7.066e-16, 7.044402e-16, 7.057663e-16, 7.015049e-16, 
    7.021938e-16, 7.017839e-16, 7.002839e-16, 7.050711e-16, 7.026159e-16, 
    7.071468e-16, 7.058192e-16, 7.096905e-16, 7.077661e-16, 7.115431e-16, 
    7.131537e-16, 7.146696e-16, 7.16437e-16, 7.014103e-16, 7.008889e-16, 
    7.018227e-16, 7.03113e-16, 7.043104e-16, 7.059002e-16, 7.060629e-16, 
    7.063604e-16, 7.071312e-16, 7.077787e-16, 7.064541e-16, 7.07941e-16, 
    7.023527e-16, 7.052842e-16, 7.006913e-16, 7.020753e-16, 7.030372e-16, 
    7.026157e-16, 7.048048e-16, 7.053201e-16, 7.074122e-16, 7.063313e-16, 
    7.12756e-16, 7.09917e-16, 7.177825e-16, 7.155886e-16, 7.007066e-16, 
    7.014087e-16, 7.038492e-16, 7.026885e-16, 7.060064e-16, 7.068218e-16, 
    7.074846e-16, 7.083309e-16, 7.084225e-16, 7.089237e-16, 7.081023e-16, 
    7.088915e-16, 7.059035e-16, 7.072396e-16, 7.035709e-16, 7.044644e-16, 
    7.040536e-16, 7.036025e-16, 7.049942e-16, 7.064748e-16, 7.065071e-16, 
    7.069814e-16, 7.08316e-16, 7.060199e-16, 7.131207e-16, 7.087384e-16, 
    7.021739e-16, 7.035238e-16, 7.037173e-16, 7.031945e-16, 7.0674e-16, 
    7.054563e-16, 7.089116e-16, 7.079787e-16, 7.095071e-16, 7.087478e-16, 
    7.08636e-16, 7.076602e-16, 7.070521e-16, 7.05515e-16, 7.042633e-16, 
    7.032704e-16, 7.035014e-16, 7.045919e-16, 7.065655e-16, 7.084306e-16, 
    7.080221e-16, 7.09391e-16, 7.057661e-16, 7.072869e-16, 7.06699e-16, 
    7.082314e-16, 7.048724e-16, 7.077312e-16, 7.041406e-16, 7.044559e-16, 
    7.054307e-16, 7.073895e-16, 7.078235e-16, 7.082855e-16, 7.080005e-16, 
    7.066157e-16, 7.063889e-16, 7.054072e-16, 7.051357e-16, 7.043873e-16, 
    7.037671e-16, 7.043336e-16, 7.049282e-16, 7.066165e-16, 7.08136e-16, 
    7.097911e-16, 7.101961e-16, 7.121253e-16, 7.105541e-16, 7.13145e-16, 
    7.109412e-16, 7.147546e-16, 7.078977e-16, 7.108777e-16, 7.054753e-16, 
    7.060584e-16, 7.071119e-16, 7.095265e-16, 7.082242e-16, 7.097475e-16, 
    7.063801e-16, 7.046292e-16, 7.041767e-16, 7.033306e-16, 7.04196e-16, 
    7.041257e-16, 7.049533e-16, 7.046874e-16, 7.066725e-16, 7.056066e-16, 
    7.08633e-16, 7.097356e-16, 7.128459e-16, 7.147487e-16, 7.166841e-16, 
    7.175373e-16, 7.17797e-16, 7.179055e-16 ;

 CWDC_TO_LITR2C =
  5.296366e-16, 5.309853e-16, 5.307233e-16, 5.3181e-16, 5.312074e-16, 
    5.319187e-16, 5.299103e-16, 5.310386e-16, 5.303186e-16, 5.297583e-16, 
    5.339154e-16, 5.318585e-16, 5.360502e-16, 5.347408e-16, 5.380277e-16, 
    5.358463e-16, 5.384671e-16, 5.379653e-16, 5.394761e-16, 5.390436e-16, 
    5.409727e-16, 5.396758e-16, 5.419722e-16, 5.406634e-16, 5.408681e-16, 
    5.396329e-16, 5.322732e-16, 5.336593e-16, 5.321909e-16, 5.323887e-16, 
    5.323001e-16, 5.312197e-16, 5.306747e-16, 5.295338e-16, 5.297411e-16, 
    5.305792e-16, 5.324776e-16, 5.318338e-16, 5.334566e-16, 5.334201e-16, 
    5.352238e-16, 5.344108e-16, 5.374386e-16, 5.36579e-16, 5.390616e-16, 
    5.384377e-16, 5.390322e-16, 5.388521e-16, 5.390346e-16, 5.381194e-16, 
    5.385116e-16, 5.377061e-16, 5.34563e-16, 5.354875e-16, 5.327278e-16, 
    5.310646e-16, 5.299598e-16, 5.291748e-16, 5.292858e-16, 5.294973e-16, 
    5.30584e-16, 5.316053e-16, 5.32383e-16, 5.329028e-16, 5.334148e-16, 
    5.349619e-16, 5.357811e-16, 5.376121e-16, 5.372823e-16, 5.378413e-16, 
    5.383757e-16, 5.392717e-16, 5.391243e-16, 5.395188e-16, 5.378269e-16, 
    5.389514e-16, 5.370943e-16, 5.376025e-16, 5.335523e-16, 5.320076e-16, 
    5.313491e-16, 5.307736e-16, 5.293711e-16, 5.303397e-16, 5.299579e-16, 
    5.308664e-16, 5.31443e-16, 5.311579e-16, 5.32917e-16, 5.322334e-16, 
    5.358295e-16, 5.342819e-16, 5.383134e-16, 5.3735e-16, 5.385442e-16, 
    5.379351e-16, 5.389784e-16, 5.380395e-16, 5.396657e-16, 5.400193e-16, 
    5.397776e-16, 5.407062e-16, 5.379874e-16, 5.390321e-16, 5.311499e-16, 
    5.311963e-16, 5.314131e-16, 5.304599e-16, 5.304017e-16, 5.29528e-16, 
    5.303056e-16, 5.306364e-16, 5.314765e-16, 5.319729e-16, 5.324446e-16, 
    5.334813e-16, 5.346376e-16, 5.362531e-16, 5.374125e-16, 5.381889e-16, 
    5.37713e-16, 5.381332e-16, 5.376634e-16, 5.374432e-16, 5.398867e-16, 
    5.385152e-16, 5.405727e-16, 5.40459e-16, 5.395281e-16, 5.404718e-16, 
    5.31229e-16, 5.309614e-16, 5.300313e-16, 5.307592e-16, 5.294328e-16, 
    5.301753e-16, 5.306018e-16, 5.322473e-16, 5.326089e-16, 5.329436e-16, 
    5.336047e-16, 5.344524e-16, 5.35938e-16, 5.372292e-16, 5.384068e-16, 
    5.383206e-16, 5.38351e-16, 5.386137e-16, 5.379625e-16, 5.387206e-16, 
    5.388476e-16, 5.385152e-16, 5.404438e-16, 5.398931e-16, 5.404566e-16, 
    5.400982e-16, 5.310484e-16, 5.314987e-16, 5.312554e-16, 5.317129e-16, 
    5.313905e-16, 5.328228e-16, 5.33252e-16, 5.352582e-16, 5.344357e-16, 
    5.35745e-16, 5.345688e-16, 5.347773e-16, 5.357869e-16, 5.346326e-16, 
    5.371577e-16, 5.354457e-16, 5.386239e-16, 5.369159e-16, 5.387308e-16, 
    5.384017e-16, 5.389467e-16, 5.394344e-16, 5.400479e-16, 5.411786e-16, 
    5.409169e-16, 5.418621e-16, 5.321699e-16, 5.327532e-16, 5.327022e-16, 
    5.333126e-16, 5.337637e-16, 5.347414e-16, 5.363073e-16, 5.357188e-16, 
    5.367993e-16, 5.37016e-16, 5.353745e-16, 5.363823e-16, 5.331437e-16, 
    5.336672e-16, 5.333558e-16, 5.322157e-16, 5.35854e-16, 5.339881e-16, 
    5.374316e-16, 5.364226e-16, 5.393648e-16, 5.379022e-16, 5.407728e-16, 
    5.419968e-16, 5.43149e-16, 5.444921e-16, 5.330718e-16, 5.326756e-16, 
    5.333853e-16, 5.343659e-16, 5.352759e-16, 5.364841e-16, 5.366078e-16, 
    5.368339e-16, 5.374197e-16, 5.379118e-16, 5.369051e-16, 5.380352e-16, 
    5.33788e-16, 5.36016e-16, 5.325254e-16, 5.335772e-16, 5.343082e-16, 
    5.339879e-16, 5.356516e-16, 5.360433e-16, 5.376333e-16, 5.368118e-16, 
    5.416946e-16, 5.395369e-16, 5.455147e-16, 5.438474e-16, 5.32537e-16, 
    5.330706e-16, 5.349254e-16, 5.340433e-16, 5.365649e-16, 5.371846e-16, 
    5.376884e-16, 5.383315e-16, 5.384011e-16, 5.38782e-16, 5.381578e-16, 
    5.387575e-16, 5.364867e-16, 5.375021e-16, 5.347139e-16, 5.35393e-16, 
    5.350807e-16, 5.347379e-16, 5.357956e-16, 5.369208e-16, 5.369454e-16, 
    5.373059e-16, 5.383202e-16, 5.365751e-16, 5.419718e-16, 5.386412e-16, 
    5.336521e-16, 5.346781e-16, 5.348251e-16, 5.344278e-16, 5.371224e-16, 
    5.361468e-16, 5.387728e-16, 5.380638e-16, 5.392254e-16, 5.386483e-16, 
    5.385633e-16, 5.378217e-16, 5.373596e-16, 5.361914e-16, 5.352401e-16, 
    5.344855e-16, 5.346611e-16, 5.354899e-16, 5.369898e-16, 5.384072e-16, 
    5.380968e-16, 5.391372e-16, 5.363822e-16, 5.37538e-16, 5.370913e-16, 
    5.382558e-16, 5.357031e-16, 5.378757e-16, 5.351468e-16, 5.353865e-16, 
    5.361274e-16, 5.37616e-16, 5.379458e-16, 5.38297e-16, 5.380804e-16, 
    5.370279e-16, 5.368556e-16, 5.361095e-16, 5.359031e-16, 5.353344e-16, 
    5.34863e-16, 5.352935e-16, 5.357454e-16, 5.370286e-16, 5.381834e-16, 
    5.394412e-16, 5.39749e-16, 5.412152e-16, 5.400211e-16, 5.419902e-16, 
    5.403153e-16, 5.432135e-16, 5.380022e-16, 5.40267e-16, 5.361613e-16, 
    5.366044e-16, 5.37405e-16, 5.392402e-16, 5.382504e-16, 5.394081e-16, 
    5.368489e-16, 5.355182e-16, 5.351743e-16, 5.345313e-16, 5.35189e-16, 
    5.351355e-16, 5.357645e-16, 5.355624e-16, 5.370711e-16, 5.36261e-16, 
    5.385611e-16, 5.393991e-16, 5.417629e-16, 5.432091e-16, 5.446799e-16, 
    5.453284e-16, 5.455257e-16, 5.456082e-16 ;

 CWDC_TO_LITR3C =
  1.672537e-16, 1.676795e-16, 1.675968e-16, 1.6794e-16, 1.677497e-16, 
    1.679743e-16, 1.673401e-16, 1.676964e-16, 1.67469e-16, 1.672921e-16, 
    1.686049e-16, 1.679553e-16, 1.69279e-16, 1.688655e-16, 1.699035e-16, 
    1.692146e-16, 1.700422e-16, 1.698838e-16, 1.703609e-16, 1.702243e-16, 
    1.708335e-16, 1.704239e-16, 1.711491e-16, 1.707358e-16, 1.708004e-16, 
    1.704104e-16, 1.680863e-16, 1.68524e-16, 1.680603e-16, 1.681228e-16, 
    1.680947e-16, 1.677536e-16, 1.675815e-16, 1.672212e-16, 1.672867e-16, 
    1.675513e-16, 1.681508e-16, 1.679475e-16, 1.6846e-16, 1.684484e-16, 
    1.69018e-16, 1.687613e-16, 1.697175e-16, 1.69446e-16, 1.7023e-16, 
    1.70033e-16, 1.702207e-16, 1.701638e-16, 1.702214e-16, 1.699325e-16, 
    1.700563e-16, 1.698019e-16, 1.688094e-16, 1.691013e-16, 1.682298e-16, 
    1.677046e-16, 1.673557e-16, 1.671078e-16, 1.671429e-16, 1.672097e-16, 
    1.675529e-16, 1.678754e-16, 1.681209e-16, 1.682851e-16, 1.684468e-16, 
    1.689353e-16, 1.69194e-16, 1.697722e-16, 1.696681e-16, 1.698446e-16, 
    1.700134e-16, 1.702963e-16, 1.702498e-16, 1.703744e-16, 1.698401e-16, 
    1.701952e-16, 1.696087e-16, 1.697692e-16, 1.684902e-16, 1.680024e-16, 
    1.677944e-16, 1.676127e-16, 1.671698e-16, 1.674757e-16, 1.673551e-16, 
    1.67642e-16, 1.678241e-16, 1.677341e-16, 1.682896e-16, 1.680737e-16, 
    1.692093e-16, 1.687206e-16, 1.699937e-16, 1.696895e-16, 1.700666e-16, 
    1.698742e-16, 1.702037e-16, 1.699072e-16, 1.704208e-16, 1.705324e-16, 
    1.704561e-16, 1.707493e-16, 1.698907e-16, 1.702207e-16, 1.677315e-16, 
    1.677462e-16, 1.678147e-16, 1.675137e-16, 1.674953e-16, 1.672194e-16, 
    1.674649e-16, 1.675694e-16, 1.678347e-16, 1.679914e-16, 1.681404e-16, 
    1.684678e-16, 1.688329e-16, 1.693431e-16, 1.697092e-16, 1.699544e-16, 
    1.698041e-16, 1.699368e-16, 1.697884e-16, 1.697189e-16, 1.704905e-16, 
    1.700574e-16, 1.707072e-16, 1.706713e-16, 1.703773e-16, 1.706753e-16, 
    1.677565e-16, 1.67672e-16, 1.673783e-16, 1.676082e-16, 1.671893e-16, 
    1.674238e-16, 1.675585e-16, 1.680781e-16, 1.681923e-16, 1.68298e-16, 
    1.685067e-16, 1.687745e-16, 1.692436e-16, 1.696513e-16, 1.700232e-16, 
    1.69996e-16, 1.700056e-16, 1.700885e-16, 1.698829e-16, 1.701223e-16, 
    1.701624e-16, 1.700574e-16, 1.706665e-16, 1.704926e-16, 1.706705e-16, 
    1.705573e-16, 1.676995e-16, 1.678417e-16, 1.677649e-16, 1.679093e-16, 
    1.678075e-16, 1.682598e-16, 1.683954e-16, 1.690289e-16, 1.687692e-16, 
    1.691826e-16, 1.688112e-16, 1.68877e-16, 1.691959e-16, 1.688313e-16, 
    1.696287e-16, 1.690881e-16, 1.700918e-16, 1.695524e-16, 1.701255e-16, 
    1.700216e-16, 1.701937e-16, 1.703477e-16, 1.705414e-16, 1.708985e-16, 
    1.708159e-16, 1.711143e-16, 1.680537e-16, 1.682379e-16, 1.682217e-16, 
    1.684145e-16, 1.68557e-16, 1.688657e-16, 1.693602e-16, 1.691744e-16, 
    1.695156e-16, 1.69584e-16, 1.690656e-16, 1.693839e-16, 1.683612e-16, 
    1.685265e-16, 1.684281e-16, 1.680681e-16, 1.692171e-16, 1.686278e-16, 
    1.697152e-16, 1.693966e-16, 1.703257e-16, 1.698639e-16, 1.707704e-16, 
    1.711569e-16, 1.715207e-16, 1.719449e-16, 1.683385e-16, 1.682133e-16, 
    1.684375e-16, 1.687471e-16, 1.690345e-16, 1.69416e-16, 1.694551e-16, 
    1.695265e-16, 1.697115e-16, 1.698669e-16, 1.69549e-16, 1.699058e-16, 
    1.685646e-16, 1.692682e-16, 1.681659e-16, 1.684981e-16, 1.687289e-16, 
    1.686278e-16, 1.691531e-16, 1.692768e-16, 1.697789e-16, 1.695195e-16, 
    1.710614e-16, 1.703801e-16, 1.722678e-16, 1.717413e-16, 1.681696e-16, 
    1.683381e-16, 1.689238e-16, 1.686453e-16, 1.694415e-16, 1.696372e-16, 
    1.697963e-16, 1.699994e-16, 1.700214e-16, 1.701417e-16, 1.699445e-16, 
    1.701339e-16, 1.694168e-16, 1.697375e-16, 1.68857e-16, 1.690715e-16, 
    1.689729e-16, 1.688646e-16, 1.691986e-16, 1.69554e-16, 1.695617e-16, 
    1.696755e-16, 1.699958e-16, 1.694448e-16, 1.71149e-16, 1.700972e-16, 
    1.685217e-16, 1.688457e-16, 1.688921e-16, 1.687667e-16, 1.696176e-16, 
    1.693095e-16, 1.701388e-16, 1.699149e-16, 1.702817e-16, 1.700995e-16, 
    1.700726e-16, 1.698384e-16, 1.696925e-16, 1.693236e-16, 1.690232e-16, 
    1.687849e-16, 1.688403e-16, 1.691021e-16, 1.695757e-16, 1.700233e-16, 
    1.699253e-16, 1.702538e-16, 1.693839e-16, 1.697488e-16, 1.696078e-16, 
    1.699755e-16, 1.691694e-16, 1.698555e-16, 1.689937e-16, 1.690694e-16, 
    1.693034e-16, 1.697735e-16, 1.698776e-16, 1.699885e-16, 1.699201e-16, 
    1.695878e-16, 1.695334e-16, 1.692977e-16, 1.692326e-16, 1.69053e-16, 
    1.689041e-16, 1.690401e-16, 1.691828e-16, 1.69588e-16, 1.699526e-16, 
    1.703499e-16, 1.704471e-16, 1.709101e-16, 1.70533e-16, 1.711548e-16, 
    1.706259e-16, 1.715411e-16, 1.698954e-16, 1.706106e-16, 1.693141e-16, 
    1.69454e-16, 1.697068e-16, 1.702864e-16, 1.699738e-16, 1.703394e-16, 
    1.695312e-16, 1.69111e-16, 1.690024e-16, 1.687994e-16, 1.69007e-16, 
    1.689902e-16, 1.691888e-16, 1.69125e-16, 1.696014e-16, 1.693456e-16, 
    1.700719e-16, 1.703366e-16, 1.71083e-16, 1.715397e-16, 1.720042e-16, 
    1.72209e-16, 1.722713e-16, 1.722973e-16 ;

 CWDC_vr =
  5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 5.110341e-05, 
    5.110342e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 
    5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110341e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 
    5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110339e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110342e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.11034e-05, 5.11034e-05, 5.110339e-05, 5.110339e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.11034e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 5.11034e-05, 
    5.110341e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.110339e-05, 
    5.110339e-05, 5.110339e-05, 5.110339e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09 ;

 CWDN_TO_LITR2N =
  1.059273e-18, 1.06197e-18, 1.061447e-18, 1.06362e-18, 1.062415e-18, 
    1.063837e-18, 1.059821e-18, 1.062077e-18, 1.060637e-18, 1.059517e-18, 
    1.067831e-18, 1.063717e-18, 1.0721e-18, 1.069482e-18, 1.076055e-18, 
    1.071693e-18, 1.076934e-18, 1.075931e-18, 1.078952e-18, 1.078087e-18, 
    1.081945e-18, 1.079351e-18, 1.083944e-18, 1.081327e-18, 1.081736e-18, 
    1.079266e-18, 1.064546e-18, 1.067319e-18, 1.064382e-18, 1.064777e-18, 
    1.0646e-18, 1.062439e-18, 1.061349e-18, 1.059067e-18, 1.059482e-18, 
    1.061158e-18, 1.064955e-18, 1.063668e-18, 1.066913e-18, 1.06684e-18, 
    1.070448e-18, 1.068822e-18, 1.074877e-18, 1.073158e-18, 1.078123e-18, 
    1.076875e-18, 1.078064e-18, 1.077704e-18, 1.078069e-18, 1.076239e-18, 
    1.077023e-18, 1.075412e-18, 1.069126e-18, 1.070975e-18, 1.065456e-18, 
    1.062129e-18, 1.05992e-18, 1.05835e-18, 1.058572e-18, 1.058995e-18, 
    1.061168e-18, 1.063211e-18, 1.064766e-18, 1.065805e-18, 1.06683e-18, 
    1.069924e-18, 1.071562e-18, 1.075224e-18, 1.074565e-18, 1.075683e-18, 
    1.076751e-18, 1.078543e-18, 1.078249e-18, 1.079038e-18, 1.075654e-18, 
    1.077903e-18, 1.074189e-18, 1.075205e-18, 1.067105e-18, 1.064015e-18, 
    1.062698e-18, 1.061547e-18, 1.058742e-18, 1.060679e-18, 1.059916e-18, 
    1.061733e-18, 1.062886e-18, 1.062316e-18, 1.065834e-18, 1.064467e-18, 
    1.071659e-18, 1.068564e-18, 1.076627e-18, 1.0747e-18, 1.077088e-18, 
    1.07587e-18, 1.077957e-18, 1.076079e-18, 1.079331e-18, 1.080039e-18, 
    1.079555e-18, 1.081412e-18, 1.075975e-18, 1.078064e-18, 1.0623e-18, 
    1.062393e-18, 1.062826e-18, 1.06092e-18, 1.060803e-18, 1.059056e-18, 
    1.060611e-18, 1.061273e-18, 1.062953e-18, 1.063946e-18, 1.064889e-18, 
    1.066962e-18, 1.069275e-18, 1.072506e-18, 1.074825e-18, 1.076378e-18, 
    1.075426e-18, 1.076266e-18, 1.075327e-18, 1.074886e-18, 1.079773e-18, 
    1.07703e-18, 1.081145e-18, 1.080918e-18, 1.079056e-18, 1.080944e-18, 
    1.062458e-18, 1.061923e-18, 1.060063e-18, 1.061519e-18, 1.058866e-18, 
    1.060351e-18, 1.061204e-18, 1.064495e-18, 1.065218e-18, 1.065887e-18, 
    1.067209e-18, 1.068905e-18, 1.071876e-18, 1.074458e-18, 1.076814e-18, 
    1.076641e-18, 1.076702e-18, 1.077227e-18, 1.075925e-18, 1.077441e-18, 
    1.077695e-18, 1.07703e-18, 1.080888e-18, 1.079786e-18, 1.080913e-18, 
    1.080196e-18, 1.062097e-18, 1.062998e-18, 1.062511e-18, 1.063426e-18, 
    1.062781e-18, 1.065646e-18, 1.066504e-18, 1.070516e-18, 1.068871e-18, 
    1.07149e-18, 1.069138e-18, 1.069555e-18, 1.071574e-18, 1.069265e-18, 
    1.074315e-18, 1.070891e-18, 1.077248e-18, 1.073832e-18, 1.077462e-18, 
    1.076803e-18, 1.077893e-18, 1.078869e-18, 1.080096e-18, 1.082357e-18, 
    1.081834e-18, 1.083724e-18, 1.06434e-18, 1.065506e-18, 1.065404e-18, 
    1.066625e-18, 1.067528e-18, 1.069483e-18, 1.072615e-18, 1.071438e-18, 
    1.073599e-18, 1.074032e-18, 1.070749e-18, 1.072765e-18, 1.066287e-18, 
    1.067335e-18, 1.066712e-18, 1.064432e-18, 1.071708e-18, 1.067976e-18, 
    1.074863e-18, 1.072845e-18, 1.07873e-18, 1.075805e-18, 1.081546e-18, 
    1.083994e-18, 1.086298e-18, 1.088984e-18, 1.066144e-18, 1.065351e-18, 
    1.06677e-18, 1.068732e-18, 1.070552e-18, 1.072968e-18, 1.073216e-18, 
    1.073668e-18, 1.074839e-18, 1.075824e-18, 1.07381e-18, 1.07607e-18, 
    1.067576e-18, 1.072032e-18, 1.065051e-18, 1.067154e-18, 1.068617e-18, 
    1.067976e-18, 1.071303e-18, 1.072087e-18, 1.075267e-18, 1.073624e-18, 
    1.083389e-18, 1.079074e-18, 1.091029e-18, 1.087695e-18, 1.065074e-18, 
    1.066141e-18, 1.069851e-18, 1.068087e-18, 1.07313e-18, 1.074369e-18, 
    1.075377e-18, 1.076663e-18, 1.076802e-18, 1.077564e-18, 1.076316e-18, 
    1.077515e-18, 1.072973e-18, 1.075004e-18, 1.069428e-18, 1.070786e-18, 
    1.070161e-18, 1.069476e-18, 1.071591e-18, 1.073842e-18, 1.073891e-18, 
    1.074612e-18, 1.07664e-18, 1.07315e-18, 1.083944e-18, 1.077282e-18, 
    1.067304e-18, 1.069356e-18, 1.06965e-18, 1.068856e-18, 1.074245e-18, 
    1.072293e-18, 1.077546e-18, 1.076128e-18, 1.078451e-18, 1.077297e-18, 
    1.077127e-18, 1.075643e-18, 1.074719e-18, 1.072383e-18, 1.07048e-18, 
    1.068971e-18, 1.069322e-18, 1.07098e-18, 1.07398e-18, 1.076814e-18, 
    1.076194e-18, 1.078274e-18, 1.072764e-18, 1.075076e-18, 1.074183e-18, 
    1.076512e-18, 1.071406e-18, 1.075751e-18, 1.070294e-18, 1.070773e-18, 
    1.072255e-18, 1.075232e-18, 1.075892e-18, 1.076594e-18, 1.076161e-18, 
    1.074056e-18, 1.073711e-18, 1.072219e-18, 1.071806e-18, 1.070669e-18, 
    1.069726e-18, 1.070587e-18, 1.071491e-18, 1.074057e-18, 1.076367e-18, 
    1.078882e-18, 1.079498e-18, 1.08243e-18, 1.080042e-18, 1.08398e-18, 
    1.080631e-18, 1.086427e-18, 1.076005e-18, 1.080534e-18, 1.072323e-18, 
    1.073209e-18, 1.07481e-18, 1.07848e-18, 1.076501e-18, 1.078816e-18, 
    1.073698e-18, 1.071036e-18, 1.070349e-18, 1.069063e-18, 1.070378e-18, 
    1.070271e-18, 1.071529e-18, 1.071125e-18, 1.074142e-18, 1.072522e-18, 
    1.077122e-18, 1.078798e-18, 1.083526e-18, 1.086418e-18, 1.08936e-18, 
    1.090657e-18, 1.091051e-18, 1.091216e-18 ;

 CWDN_TO_LITR3N =
  3.345073e-19, 3.353591e-19, 3.351936e-19, 3.3588e-19, 3.354994e-19, 
    3.359487e-19, 3.346802e-19, 3.353928e-19, 3.34938e-19, 3.345842e-19, 
    3.372097e-19, 3.359106e-19, 3.38558e-19, 3.377311e-19, 3.39807e-19, 
    3.384292e-19, 3.400845e-19, 3.397676e-19, 3.407218e-19, 3.404486e-19, 
    3.41667e-19, 3.408479e-19, 3.422982e-19, 3.414716e-19, 3.416009e-19, 
    3.408208e-19, 3.361725e-19, 3.37048e-19, 3.361206e-19, 3.362455e-19, 
    3.361895e-19, 3.355072e-19, 3.351629e-19, 3.344424e-19, 3.345733e-19, 
    3.351026e-19, 3.363017e-19, 3.358951e-19, 3.3692e-19, 3.368969e-19, 
    3.380361e-19, 3.375226e-19, 3.394349e-19, 3.38892e-19, 3.4046e-19, 
    3.400659e-19, 3.404414e-19, 3.403276e-19, 3.404429e-19, 3.398649e-19, 
    3.401126e-19, 3.396039e-19, 3.376188e-19, 3.382026e-19, 3.364597e-19, 
    3.354092e-19, 3.347114e-19, 3.342157e-19, 3.342858e-19, 3.344193e-19, 
    3.351057e-19, 3.357507e-19, 3.362419e-19, 3.365702e-19, 3.368935e-19, 
    3.378707e-19, 3.38388e-19, 3.395445e-19, 3.393362e-19, 3.396892e-19, 
    3.400267e-19, 3.405926e-19, 3.404996e-19, 3.407487e-19, 3.396801e-19, 
    3.403904e-19, 3.392174e-19, 3.395384e-19, 3.369804e-19, 3.360048e-19, 
    3.355889e-19, 3.352254e-19, 3.343396e-19, 3.349514e-19, 3.347103e-19, 
    3.35284e-19, 3.356482e-19, 3.354681e-19, 3.365791e-19, 3.361474e-19, 
    3.384187e-19, 3.374412e-19, 3.399874e-19, 3.39379e-19, 3.401332e-19, 
    3.397485e-19, 3.404074e-19, 3.398144e-19, 3.408415e-19, 3.410648e-19, 
    3.409122e-19, 3.414986e-19, 3.397815e-19, 3.404413e-19, 3.35463e-19, 
    3.354924e-19, 3.356293e-19, 3.350273e-19, 3.349905e-19, 3.344387e-19, 
    3.349299e-19, 3.351388e-19, 3.356694e-19, 3.359829e-19, 3.362808e-19, 
    3.369355e-19, 3.376658e-19, 3.386861e-19, 3.394184e-19, 3.399088e-19, 
    3.396082e-19, 3.398736e-19, 3.395769e-19, 3.394378e-19, 3.409811e-19, 
    3.401149e-19, 3.414143e-19, 3.413425e-19, 3.407546e-19, 3.413506e-19, 
    3.355131e-19, 3.35344e-19, 3.347566e-19, 3.352164e-19, 3.343786e-19, 
    3.348475e-19, 3.351169e-19, 3.361562e-19, 3.363846e-19, 3.365959e-19, 
    3.370135e-19, 3.375489e-19, 3.384871e-19, 3.393026e-19, 3.400464e-19, 
    3.39992e-19, 3.400111e-19, 3.401771e-19, 3.397658e-19, 3.402446e-19, 
    3.403248e-19, 3.401149e-19, 3.413329e-19, 3.409851e-19, 3.41341e-19, 
    3.411146e-19, 3.35399e-19, 3.356834e-19, 3.355297e-19, 3.358186e-19, 
    3.35615e-19, 3.365197e-19, 3.367907e-19, 3.380578e-19, 3.375383e-19, 
    3.383652e-19, 3.376225e-19, 3.377541e-19, 3.383918e-19, 3.376627e-19, 
    3.392575e-19, 3.381762e-19, 3.401835e-19, 3.391048e-19, 3.40251e-19, 
    3.400432e-19, 3.403874e-19, 3.406954e-19, 3.410829e-19, 3.41797e-19, 
    3.416317e-19, 3.422287e-19, 3.361073e-19, 3.364757e-19, 3.364435e-19, 
    3.36829e-19, 3.371139e-19, 3.377314e-19, 3.387204e-19, 3.383487e-19, 
    3.390311e-19, 3.39168e-19, 3.381313e-19, 3.387678e-19, 3.367224e-19, 
    3.37053e-19, 3.368563e-19, 3.361363e-19, 3.384341e-19, 3.372556e-19, 
    3.394305e-19, 3.387932e-19, 3.406515e-19, 3.397277e-19, 3.415407e-19, 
    3.423138e-19, 3.430414e-19, 3.438897e-19, 3.366769e-19, 3.364267e-19, 
    3.368749e-19, 3.374942e-19, 3.38069e-19, 3.388321e-19, 3.389102e-19, 
    3.39053e-19, 3.39423e-19, 3.397338e-19, 3.390979e-19, 3.398117e-19, 
    3.371293e-19, 3.385364e-19, 3.363318e-19, 3.369961e-19, 3.374578e-19, 
    3.372555e-19, 3.383063e-19, 3.385537e-19, 3.395578e-19, 3.39039e-19, 
    3.421229e-19, 3.407602e-19, 3.445356e-19, 3.434825e-19, 3.363392e-19, 
    3.366762e-19, 3.378476e-19, 3.372905e-19, 3.388831e-19, 3.392745e-19, 
    3.395926e-19, 3.399988e-19, 3.400428e-19, 3.402834e-19, 3.398891e-19, 
    3.402679e-19, 3.388337e-19, 3.39475e-19, 3.37714e-19, 3.381429e-19, 
    3.379457e-19, 3.377292e-19, 3.383972e-19, 3.391079e-19, 3.391234e-19, 
    3.393511e-19, 3.399917e-19, 3.388895e-19, 3.42298e-19, 3.401944e-19, 
    3.370435e-19, 3.376914e-19, 3.377843e-19, 3.375333e-19, 3.392352e-19, 
    3.38619e-19, 3.402776e-19, 3.398298e-19, 3.405634e-19, 3.401989e-19, 
    3.401452e-19, 3.396769e-19, 3.39385e-19, 3.386472e-19, 3.380464e-19, 
    3.375698e-19, 3.376807e-19, 3.382041e-19, 3.391514e-19, 3.400467e-19, 
    3.398506e-19, 3.405077e-19, 3.387677e-19, 3.394977e-19, 3.392155e-19, 
    3.39951e-19, 3.383388e-19, 3.39711e-19, 3.379875e-19, 3.381388e-19, 
    3.386068e-19, 3.395469e-19, 3.397553e-19, 3.39977e-19, 3.398403e-19, 
    3.391755e-19, 3.390667e-19, 3.385955e-19, 3.384651e-19, 3.381059e-19, 
    3.378082e-19, 3.380801e-19, 3.383655e-19, 3.391759e-19, 3.399053e-19, 
    3.406997e-19, 3.408941e-19, 3.418201e-19, 3.41066e-19, 3.423096e-19, 
    3.412518e-19, 3.430822e-19, 3.397909e-19, 3.412213e-19, 3.386281e-19, 
    3.38908e-19, 3.394137e-19, 3.405727e-19, 3.399476e-19, 3.406788e-19, 
    3.390625e-19, 3.38222e-19, 3.380048e-19, 3.375987e-19, 3.380141e-19, 
    3.379803e-19, 3.383776e-19, 3.3825e-19, 3.392028e-19, 3.386912e-19, 
    3.401438e-19, 3.406731e-19, 3.42166e-19, 3.430794e-19, 3.440084e-19, 
    3.444179e-19, 3.445426e-19, 3.445946e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  2.413656e-36, 2.065401e-35, 1.367197e-35, 7.458777e-35, 2.924233e-35, 
    8.819833e-35, 3.748208e-36, 2.246482e-35, 7.197595e-36, 2.935293e-36, 
    1.796957e-33, 8.037766e-35, 3.922441e-32, 6.007093e-33, 6.052333e-31, 
    2.939911e-32, 1.094422e-30, 5.556852e-31, 4.175555e-30, 2.359349e-30, 
    2.893847e-29, 5.424175e-30, 1.017046e-28, 1.948533e-29, 2.531664e-29, 
    5.128552e-30, 1.5186e-34, 1.229759e-33, 1.339012e-34, 1.812237e-34, 
    1.582295e-34, 2.981927e-35, 1.267358e-35, 2.04289e-36, 2.854736e-36, 
    1.088977e-35, 2.075535e-34, 7.733206e-35, 9.06774e-34, 8.585492e-34, 
    1.206895e-32, 3.712564e-33, 2.708682e-31, 8.236855e-32, 2.416494e-30, 
    1.051322e-30, 2.324528e-30, 1.82943e-30, 2.331775e-30, 6.847458e-31, 
    1.161084e-30, 3.905416e-31, 4.637344e-33, 1.761981e-32, 3.033677e-34, 
    2.342121e-35, 4.05827e-36, 1.140883e-36, 1.366814e-36, 1.926661e-36, 
    1.097471e-35, 5.431533e-35, 1.795261e-34, 3.950291e-34, 8.518304e-34, 
    8.288211e-33, 2.678748e-32, 3.436761e-31, 2.184636e-31, 4.697071e-31, 
    9.671604e-31, 3.190841e-30, 2.625917e-30, 4.41738e-30, 4.603185e-31, 
    2.088884e-30, 1.685259e-31, 3.389846e-31, 1.048926e-33, 1.010662e-34, 
    3.652738e-35, 1.480341e-35, 1.570089e-36, 7.446789e-36, 4.047018e-36, 
    1.712407e-35, 4.221452e-35, 2.705511e-35, 4.035902e-34, 1.42863e-34, 
    2.869719e-32, 3.075397e-33, 8.894096e-31, 2.398156e-31, 1.212633e-30, 
    5.331979e-31, 2.164703e-30, 6.143018e-31, 5.354316e-30, 8.491746e-30, 
    6.198718e-30, 2.057202e-29, 5.724397e-31, 2.324658e-30, 2.671984e-35, 
    2.873639e-35, 4.028986e-35, 9.014748e-36, 8.217192e-36, 2.024267e-36, 
    7.050135e-36, 1.192036e-35, 4.446345e-35, 9.581258e-35, 1.972759e-34, 
    9.40965e-34, 5.171452e-33, 5.218879e-32, 2.613056e-31, 7.518973e-31, 
    3.941118e-31, 6.973537e-31, 3.683514e-31, 2.724792e-31, 7.147453e-30, 
    1.166841e-30, 1.73386e-29, 1.498157e-29, 4.472238e-30, 1.523048e-29, 
    3.024102e-35, 1.988205e-35, 4.550449e-36, 1.44646e-35, 1.73507e-36, 
    5.729078e-36, 1.12904e-35, 1.460426e-34, 2.53197e-34, 4.202358e-34, 
    1.130701e-33, 3.94548e-33, 3.344858e-32, 2.031258e-31, 1.00837e-30, 
    8.979328e-31, 9.353917e-31, 1.33104e-30, 5.534872e-31, 1.535411e-30, 
    1.819247e-30, 1.166494e-30, 1.469084e-29, 7.203947e-30, 1.493503e-29, 
    9.401376e-30, 2.279148e-35, 4.603192e-35, 3.151121e-35, 6.416304e-35, 
    3.891003e-35, 3.504587e-34, 6.685744e-34, 1.269163e-32, 3.850616e-33, 
    2.54377e-32, 4.67595e-33, 6.33306e-33, 2.703684e-32, 5.129652e-33, 
    1.84164e-31, 1.661233e-32, 1.349351e-30, 1.31887e-31, 1.556519e-30, 
    1.001499e-30, 2.074591e-30, 3.953509e-30, 8.809192e-30, 3.754736e-29, 
    2.692728e-29, 8.862534e-29, 1.296324e-34, 3.153121e-34, 2.916695e-34, 
    7.313115e-34, 1.432144e-33, 6.009421e-33, 5.630612e-32, 2.449265e-32, 
    1.119704e-31, 1.512694e-31, 1.497909e-32, 6.257924e-32, 5.680003e-34, 
    1.242106e-33, 7.802933e-34, 1.391165e-34, 2.970523e-32, 1.996976e-33, 
    2.682689e-31, 6.618635e-32, 3.607827e-30, 5.103762e-31, 2.240553e-29, 
    1.049413e-28, 4.315611e-28, 2.151595e-27, 5.097033e-34, 2.801228e-34, 
    8.151042e-34, 3.479038e-33, 1.300711e-32, 7.215027e-32, 8.574919e-32, 
    1.175121e-31, 2.638394e-31, 5.166526e-31, 1.297972e-31, 6.107406e-31, 
    1.487772e-33, 3.735418e-32, 2.231189e-34, 1.086605e-33, 3.196354e-33, 
    1.995071e-33, 2.225378e-32, 3.879716e-32, 3.537037e-31, 1.139286e-31, 
    7.1979e-29, 4.527107e-30, 7.072285e-27, 1.001204e-27, 2.26989e-34, 
    5.086269e-34, 7.850772e-33, 2.164587e-33, 8.075713e-32, 1.909646e-31, 
    3.810726e-31, 9.116114e-31, 1.000794e-30, 1.666826e-30, 7.208881e-31, 
    1.612822e-30, 7.241077e-32, 2.954449e-31, 5.773067e-33, 1.538488e-32, 
    9.818068e-33, 5.978102e-33, 2.731482e-32, 1.326861e-31, 1.371577e-31, 
    2.257592e-31, 9.004322e-31, 8.191729e-32, 1.019036e-28, 1.384652e-30, 
    1.213156e-33, 5.487309e-33, 6.787049e-33, 3.804815e-33, 1.752723e-31, 
    4.491113e-32, 1.646268e-30, 6.348694e-31, 3.001185e-30, 1.393988e-30, 
    1.244232e-30, 4.570806e-31, 2.430007e-31, 4.783712e-32, 1.235653e-32, 
    4.139165e-33, 5.346258e-33, 1.767639e-32, 1.459641e-31, 1.009369e-30, 
    6.642821e-31, 2.670752e-30, 6.253374e-32, 3.104628e-31, 1.679492e-31, 
    8.230366e-31, 2.39545e-32, 4.932957e-31, 1.079973e-32, 1.5238e-32, 
    4.370052e-32, 3.45641e-31, 5.410543e-31, 8.702187e-31, 6.493018e-31, 
    1.538556e-31, 1.211231e-31, 4.260206e-32, 3.183188e-32, 1.413956e-32, 
    7.167403e-33, 1.333833e-32, 2.544929e-32, 1.539362e-31, 7.466343e-31, 
    3.989861e-30, 5.969769e-30, 3.938643e-29, 8.521178e-30, 1.042838e-28, 
    1.24947e-29, 4.677264e-28, 5.850539e-31, 1.171975e-29, 4.582477e-32, 
    8.533778e-32, 2.588349e-31, 3.063866e-30, 8.169875e-31, 3.821891e-30, 
    1.199891e-31, 1.841584e-32, 1.123526e-32, 4.426199e-33, 1.147535e-32, 
    1.062511e-32, 2.613189e-32, 1.959549e-32, 1.632738e-31, 5.273784e-32, 
    1.240751e-30, 3.776026e-30, 7.832231e-29, 4.6458e-28, 2.680098e-27, 
    5.702732e-27, 7.160027e-27, 7.872312e-27 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  7.623649e-08, 7.644516e-08, 7.640461e-08, 7.657286e-08, 7.647954e-08, 
    7.658971e-08, 7.627882e-08, 7.645342e-08, 7.634197e-08, 7.62553e-08, 
    7.689925e-08, 7.658038e-08, 7.723048e-08, 7.70272e-08, 7.753781e-08, 
    7.719884e-08, 7.760615e-08, 7.752807e-08, 7.776314e-08, 7.76958e-08, 
    7.799632e-08, 7.779421e-08, 7.815211e-08, 7.794808e-08, 7.797998e-08, 
    7.778754e-08, 7.664459e-08, 7.685954e-08, 7.663184e-08, 7.66625e-08, 
    7.664875e-08, 7.648146e-08, 7.639712e-08, 7.622056e-08, 7.625263e-08, 
    7.638231e-08, 7.667629e-08, 7.657653e-08, 7.682798e-08, 7.682231e-08, 
    7.710213e-08, 7.697598e-08, 7.744618e-08, 7.731258e-08, 7.769862e-08, 
    7.760154e-08, 7.769405e-08, 7.766601e-08, 7.769442e-08, 7.755205e-08, 
    7.761304e-08, 7.748777e-08, 7.69996e-08, 7.714308e-08, 7.671504e-08, 
    7.64575e-08, 7.628647e-08, 7.616506e-08, 7.618222e-08, 7.621494e-08, 
    7.638307e-08, 7.654115e-08, 7.666159e-08, 7.674213e-08, 7.682149e-08, 
    7.706157e-08, 7.718869e-08, 7.747317e-08, 7.742187e-08, 7.750881e-08, 
    7.759189e-08, 7.773131e-08, 7.770838e-08, 7.776979e-08, 7.750653e-08, 
    7.768149e-08, 7.739264e-08, 7.747165e-08, 7.684295e-08, 7.660345e-08, 
    7.650154e-08, 7.64124e-08, 7.619542e-08, 7.634526e-08, 7.628619e-08, 
    7.642673e-08, 7.651601e-08, 7.647186e-08, 7.674434e-08, 7.663841e-08, 
    7.719622e-08, 7.695601e-08, 7.758219e-08, 7.74324e-08, 7.76181e-08, 
    7.752336e-08, 7.768568e-08, 7.75396e-08, 7.779266e-08, 7.784774e-08, 
    7.781009e-08, 7.795472e-08, 7.753149e-08, 7.769404e-08, 7.647062e-08, 
    7.647782e-08, 7.651137e-08, 7.636387e-08, 7.635484e-08, 7.621968e-08, 
    7.633997e-08, 7.639117e-08, 7.65212e-08, 7.659807e-08, 7.667116e-08, 
    7.683181e-08, 7.701119e-08, 7.726197e-08, 7.744212e-08, 7.756284e-08, 
    7.748882e-08, 7.755416e-08, 7.748111e-08, 7.744688e-08, 7.782709e-08, 
    7.761361e-08, 7.793392e-08, 7.791621e-08, 7.777125e-08, 7.791819e-08, 
    7.648288e-08, 7.644144e-08, 7.629752e-08, 7.641015e-08, 7.620496e-08, 
    7.631981e-08, 7.638584e-08, 7.66406e-08, 7.669659e-08, 7.674847e-08, 
    7.685095e-08, 7.698243e-08, 7.721304e-08, 7.741363e-08, 7.759672e-08, 
    7.758331e-08, 7.758803e-08, 7.762892e-08, 7.752763e-08, 7.764555e-08, 
    7.766533e-08, 7.76136e-08, 7.791383e-08, 7.782807e-08, 7.791583e-08, 
    7.785999e-08, 7.645492e-08, 7.652464e-08, 7.648696e-08, 7.65578e-08, 
    7.650789e-08, 7.672979e-08, 7.679631e-08, 7.710752e-08, 7.697984e-08, 
    7.718307e-08, 7.700049e-08, 7.703284e-08, 7.718965e-08, 7.701037e-08, 
    7.740255e-08, 7.713665e-08, 7.76305e-08, 7.736501e-08, 7.764714e-08, 
    7.759594e-08, 7.768072e-08, 7.775665e-08, 7.785217e-08, 7.802836e-08, 
    7.798757e-08, 7.813491e-08, 7.662858e-08, 7.671898e-08, 7.671105e-08, 
    7.680566e-08, 7.687562e-08, 7.702726e-08, 7.727039e-08, 7.717897e-08, 
    7.73468e-08, 7.738048e-08, 7.712552e-08, 7.728205e-08, 7.67795e-08, 
    7.686069e-08, 7.681236e-08, 7.66357e-08, 7.720001e-08, 7.691045e-08, 
    7.744509e-08, 7.728828e-08, 7.774582e-08, 7.751829e-08, 7.796511e-08, 
    7.815598e-08, 7.833569e-08, 7.854553e-08, 7.676834e-08, 7.670692e-08, 
    7.681692e-08, 7.696904e-08, 7.711023e-08, 7.729785e-08, 7.731705e-08, 
    7.735219e-08, 7.744323e-08, 7.751974e-08, 7.736328e-08, 7.753892e-08, 
    7.687949e-08, 7.722515e-08, 7.668368e-08, 7.684673e-08, 7.696008e-08, 
    7.691038e-08, 7.716854e-08, 7.722935e-08, 7.747646e-08, 7.734874e-08, 
    7.810886e-08, 7.777265e-08, 7.870533e-08, 7.844478e-08, 7.668545e-08, 
    7.676814e-08, 7.705584e-08, 7.691897e-08, 7.731038e-08, 7.740669e-08, 
    7.748498e-08, 7.758503e-08, 7.759585e-08, 7.765512e-08, 7.755798e-08, 
    7.765129e-08, 7.729825e-08, 7.745604e-08, 7.702298e-08, 7.71284e-08, 
    7.707991e-08, 7.702671e-08, 7.71909e-08, 7.736573e-08, 7.736951e-08, 
    7.742555e-08, 7.758342e-08, 7.731197e-08, 7.815218e-08, 7.763335e-08, 
    7.68583e-08, 7.701748e-08, 7.704026e-08, 7.697859e-08, 7.739703e-08, 
    7.724544e-08, 7.765367e-08, 7.754338e-08, 7.77241e-08, 7.76343e-08, 
    7.762108e-08, 7.750573e-08, 7.74339e-08, 7.725239e-08, 7.710467e-08, 
    7.698755e-08, 7.701478e-08, 7.714345e-08, 7.737644e-08, 7.759681e-08, 
    7.754854e-08, 7.771037e-08, 7.728201e-08, 7.746164e-08, 7.739221e-08, 
    7.757325e-08, 7.717654e-08, 7.751427e-08, 7.709018e-08, 7.712737e-08, 
    7.724243e-08, 7.74738e-08, 7.752503e-08, 7.757966e-08, 7.754596e-08, 
    7.738236e-08, 7.735557e-08, 7.723964e-08, 7.720762e-08, 7.711928e-08, 
    7.704612e-08, 7.711296e-08, 7.718313e-08, 7.738244e-08, 7.7562e-08, 
    7.775772e-08, 7.780563e-08, 7.803415e-08, 7.784809e-08, 7.815506e-08, 
    7.789401e-08, 7.834588e-08, 7.753389e-08, 7.788639e-08, 7.724768e-08, 
    7.731652e-08, 7.744099e-08, 7.772646e-08, 7.757239e-08, 7.775259e-08, 
    7.735452e-08, 7.714787e-08, 7.709443e-08, 7.699466e-08, 7.709671e-08, 
    7.708842e-08, 7.718606e-08, 7.715469e-08, 7.738906e-08, 7.726317e-08, 
    7.762075e-08, 7.775118e-08, 7.811946e-08, 7.834512e-08, 7.857481e-08, 
    7.867618e-08, 7.870703e-08, 7.871993e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -1.351779e-14, -1.49097e-14, -1.486075e-14, -5.998742e-15, -1.424264e-14, 
    -1.076638e-14, -2.159773e-14, -1.398267e-14, -1.559314e-14, 
    -1.507395e-14, -9.89055e-15, -1.807352e-14, -9.384968e-15, -1.067309e-14, 
    -1.464065e-14, -9.392316e-15, -1.122709e-14, -1.999415e-14, 
    -6.334882e-15, -7.596656e-15, -1.103094e-14, -1.012839e-14, 
    -1.634444e-14, -9.276045e-15, -3.617183e-15, -1.955617e-14, 
    -1.041116e-14, -8.936573e-15, -7.399145e-15, -1.231595e-14, 
    -4.472331e-15, -1.0991e-14, -1.542129e-14, -1.594805e-15, -1.922421e-14, 
    -7.5159e-15, -1.28132e-14, -1.166699e-14, -1.096666e-14, -1.729714e-14, 
    -1.644735e-14, -1.254516e-14, -1.125768e-14, -1.421534e-14, 
    -8.326944e-15, -1.418321e-14, -2.143206e-14, -9.337202e-15, 
    -6.936928e-15, -2.099415e-14, -1.545682e-14, -1.547641e-14, 
    -1.254214e-14, -1.107779e-14, -8.004355e-15, -1.386787e-16, 
    -1.127309e-14, -2.316826e-14, -1.68619e-14, -9.359954e-15, -1.37685e-14, 
    -1.910438e-14, -1.501813e-14, -1.736436e-14, -1.77797e-14, -1.319611e-14, 
    -1.586161e-14, -1.538899e-14, -1.116563e-14, -9.534187e-15, 
    -1.397136e-14, -1.138373e-14, -2.119491e-14, -1.363583e-14, -1.1369e-14, 
    -8.626683e-15, -6.13519e-15, -1.218179e-14, -1.323291e-14, -1.65882e-14, 
    -1.319153e-14, -1.410344e-14, -2.058893e-14, -1.804452e-15, 
    -1.257088e-14, -8.128182e-15, -1.044895e-14, -1.811099e-14, 
    -1.200356e-14, -1.022521e-14, -2.021431e-14, -6.981792e-15, 
    -2.056909e-14, -1.324394e-14, -1.100699e-14, -1.029181e-14, 
    -1.846813e-14, -8.294553e-15, -6.813446e-15, -7.744774e-15, 
    -7.737928e-15, -1.340767e-14, -1.609357e-14, -1.728318e-14, 
    -1.068034e-14, -9.154306e-15, -2.340413e-14, -1.852776e-14, 
    -1.370586e-14, -1.217431e-14, -1.326122e-14, -1.298369e-14, 
    -1.585637e-14, -1.57981e-14, -7.10625e-15, -6.903745e-15, -1.483808e-14, 
    -1.870938e-14, -1.223004e-14, -1.497722e-14, -1.622536e-14, 
    -9.738774e-15, -1.460767e-14, -1.258851e-14, -1.393124e-14, 
    -1.559372e-14, -1.132698e-14, -1.00458e-14, -1.720481e-14, -1.507371e-14, 
    -1.825464e-14, -1.856336e-14, -9.959086e-15, -1.031986e-14, 
    -8.840719e-15, -1.158547e-14, -8.142366e-15, -1.541591e-14, 
    -1.621065e-14, -1.175465e-14, -6.398233e-15, -1.667906e-14, 
    -1.124805e-14, -1.124329e-14, -1.40911e-14, -1.440609e-14, -1.187022e-14, 
    -7.436991e-15, -1.978893e-14, -1.692911e-14, -1.248005e-14, 
    -8.109633e-15, -1.192523e-14, -1.469813e-14, -1.421613e-14, 
    -9.133581e-15, -1.48595e-14, -1.343653e-14, -1.982535e-14, -2.161525e-14, 
    -1.407301e-14, -1.321393e-14, -4.777705e-15, -1.206904e-14, 
    -5.232109e-15, -8.490431e-15, -8.296189e-15, -1.137253e-14, 
    -1.203506e-14, -1.222937e-14, -1.564501e-14, -1.370843e-14, 
    -1.673356e-14, -1.903859e-14, -1.674877e-14, -1.477117e-14, 
    -1.170971e-14, -2.170247e-14, -1.295776e-14, -1.830823e-14, 
    -1.033203e-14, -1.562713e-14, -1.506758e-14, -9.161084e-15, 
    -1.142183e-14, -1.567202e-14, -1.135635e-14, -5.642509e-15, 
    -1.467577e-14, 2.765047e-15, -1.189569e-14, -1.591639e-14, -5.765798e-15, 
    -1.483146e-14, -1.275517e-14, -5.774497e-15, -1.154548e-14, 
    -1.587918e-14, -1.112904e-14, -5.58361e-15, -4.242229e-15, -1.02732e-14, 
    -1.848576e-14, -1.226282e-14, -1.220676e-14, -8.807383e-15, -1.83613e-14, 
    -1.28388e-14, -9.920932e-15, -2.319301e-14, -1.109264e-14, -1.425745e-14, 
    -1.447275e-14, -7.962733e-15, -1.66353e-14, -5.963053e-15, -1.674108e-14, 
    -1.120968e-14, -9.417341e-15, -1.300874e-14, -3.247895e-15, 
    -1.500845e-14, -1.92475e-14, -1.872047e-14, -1.795078e-14, -5.935256e-15, 
    -1.784417e-14, -1.271263e-14, -1.626132e-14, -9.194417e-15, 
    -1.164001e-14, -1.222978e-14, -1.367916e-14, -2.189358e-15, 
    -1.627227e-14, -1.278858e-14, -1.638685e-14, -1.039414e-14, 
    -1.197293e-14, -1.351743e-14, -9.169187e-15, -9.056902e-15, -1.12853e-14, 
    -9.347432e-15, -5.567454e-15, -2.115307e-14, -4.653202e-15, 
    -1.594008e-14, -1.352236e-14, -1.299641e-14, -1.16666e-14, -1.440868e-14, 
    -7.345354e-15, -1.641458e-14, -6.977186e-15, -7.663099e-15, -1.64278e-14, 
    -1.877748e-14, -1.32887e-14, -1.711593e-14, -1.615664e-14, -1.298796e-14, 
    -1.625307e-14, -8.719207e-15, -1.504383e-14, -1.184954e-14, 
    -7.458307e-15, -2.396503e-14, -9.46395e-15, -9.304528e-15, -9.940629e-15, 
    -1.180415e-14, -1.251617e-14, -1.368224e-14, -1.409344e-14, 
    -1.661055e-14, -1.208305e-14, -1.602872e-14, -1.696098e-14, 
    -1.553794e-15, -1.710137e-14, -1.614977e-14, -1.773117e-14, 
    -1.272687e-14, -8.183518e-15, -1.558919e-14, -1.057458e-14, -1.53328e-14, 
    -1.566878e-14, -1.439931e-14, -9.075549e-15, -1.670609e-14, 
    -1.200256e-14, -1.533652e-14, -1.050422e-14, -2.219152e-14, 
    -1.093384e-14, -1.412622e-14, -7.84617e-15, -1.050905e-14, -1.990321e-14, 
    -1.377649e-14, -1.616831e-14, -1.416724e-14, -2.013573e-14, -8.62897e-15, 
    -1.445235e-14, -1.006297e-14, -1.339319e-14, -2.047502e-14, 
    -1.196347e-14, -8.767508e-15, -1.276578e-14, -1.198794e-14, 
    -1.629174e-14, -1.701643e-14, -1.018044e-14, -1.359301e-14, 
    -1.211291e-14, -1.025095e-14, -1.139754e-14, -5.271434e-15, -1.34976e-14, 
    -1.454699e-14, -1.458996e-14, -1.634646e-14, -1.698104e-14, 
    -1.067557e-14, -1.809163e-14, -1.435599e-14, -1.00964e-14, -9.520488e-15, 
    -1.107725e-14, -1.602572e-14, -1.257202e-15, -7.90552e-15, -1.024937e-14, 
    -1.441601e-14 ;

 ERRSOI =
  -4.238846e-10, -2.284053e-10, -1.591455e-10, -3.289363e-10, -1.689234e-10, 
    -1.587468e-10, -9.051422e-11, -2.436741e-11, -4.201903e-11, 
    -2.946826e-10, -1.82126e-10, -1.574261e-10, -3.644364e-10, -4.107814e-10, 
    -3.533081e-10, -6.03723e-10, -3.862379e-10, -4.640381e-10, -2.527313e-10, 
    -3.514631e-10, -3.674683e-10, -1.452741e-10, -1.677888e-10, 
    -4.071468e-10, -2.953527e-10, -4.059214e-10, -1.85454e-10, -2.134034e-10, 
    -1.711785e-10, 3.061442e-12, -2.943318e-10, -3.392404e-10, -2.112934e-10, 
    -3.775051e-10, -3.258407e-10, -2.282697e-10, -2.68993e-10, -1.393429e-10, 
    -2.654544e-10, -4.017215e-10, -4.011136e-10, -3.907843e-10, 
    -3.184037e-10, -4.491018e-10, -3.563105e-10, -4.065293e-10, 
    -2.416013e-10, -4.400514e-10, -3.33485e-10, -2.181149e-10, -4.172998e-10, 
    -4.097254e-10, -2.912051e-10, -2.695367e-10, -4.646594e-10, 
    -2.092466e-10, -1.868514e-10, -4.066839e-10, -4.227034e-10, 
    -2.091077e-10, -3.765286e-10, -2.636567e-10, -2.66949e-10, -3.43256e-11, 
    -2.917669e-10, -2.077207e-10, -3.582299e-10, -6.747917e-10, 
    -3.667893e-10, -1.989398e-10, -2.810488e-10, -2.624057e-10, 
    -1.250253e-10, -3.205502e-10, -5.304152e-10, -3.536475e-10, -3.16265e-10, 
    -2.846573e-10, -2.316882e-10, -2.715445e-10, -2.092144e-10, 
    -3.463553e-10, -3.874743e-10, -2.307129e-10, -2.844394e-10, 
    -2.799255e-10, -9.62191e-11, -9.04289e-11, -4.91978e-10, -8.233092e-11, 
    -4.503152e-10, -9.160379e-11, -3.174412e-10, -4.001061e-10, 
    -6.737079e-10, -5.361679e-10, -3.470357e-10, -3.983806e-10, 
    -3.841449e-10, -3.944344e-10, -4.02445e-10, -1.713367e-10, -2.048916e-10, 
    -3.127986e-10, -3.314813e-10, -4.516752e-10, -2.110972e-10, 
    -4.298897e-10, -7.866774e-11, -3.993159e-10, -2.751454e-10, 
    -1.321956e-10, -1.938466e-10, -2.390089e-10, -3.28163e-10, -2.016725e-10, 
    -5.72192e-10, -2.787316e-10, -3.165934e-10, -2.85772e-10, -2.559306e-10, 
    -3.135638e-10, -4.27965e-10, -2.988979e-10, -5.375831e-10, -6.726845e-10, 
    -1.630698e-10, -1.097666e-10, -2.749034e-10, -3.680595e-10, 
    -4.244864e-10, -3.681588e-10, -1.677673e-10, -3.041394e-10, 
    -1.406784e-10, -3.4143e-10, -2.650913e-10, -2.295332e-10, -1.105021e-10, 
    -2.737246e-10, -3.96368e-10, -1.907761e-10, -3.619488e-10, -3.343566e-10, 
    -2.598341e-10, -2.177126e-10, -4.11202e-10, -5.229492e-10, -4.350253e-10, 
    -3.165385e-10, -3.66016e-10, -4.017567e-10, -1.690451e-10, -3.661287e-10, 
    -1.26777e-10, -3.363841e-10, -4.072363e-10, -1.274762e-10, -1.490979e-10, 
    5.746005e-11, -2.405864e-10, -2.613815e-10, -1.303497e-10, -2.641232e-10, 
    -1.348385e-10, -4.9125e-10, -4.067237e-10, -2.586877e-10, -3.99642e-10, 
    -3.511838e-10, -3.045844e-10, -3.24224e-10, -2.534169e-10, -3.468642e-10, 
    -3.632854e-10, -4.143118e-10, -2.629435e-10, -2.44824e-10, -3.573147e-10, 
    -4.570626e-10, -4.219037e-10, -5.191911e-10, -1.84436e-10, -3.485237e-10, 
    -1.814241e-10, -2.397006e-10, -3.837156e-10, -3.854592e-10, 
    -5.120259e-10, -2.86455e-10, -3.783383e-10, -2.117628e-10, -5.054982e-10, 
    -3.325508e-10, -1.8808e-10, -3.074666e-10, -3.586975e-10, -4.470127e-10, 
    -4.828297e-10, -3.03389e-10, -2.413825e-10, -4.818076e-10, -2.245375e-10, 
    -4.62194e-10, -1.755673e-10, -3.523277e-10, -2.846782e-10, -8.087948e-11, 
    -2.424517e-10, -2.573613e-10, -2.575671e-10, -4.206752e-10, 
    -4.151733e-10, -4.912686e-10, -2.612125e-10, -4.854672e-10, 
    -4.627518e-10, -3.674352e-10, -4.350492e-10, -4.122281e-10, 
    -2.478382e-10, -3.946881e-10, -1.149049e-10, -3.962779e-10, 
    -3.184141e-10, -3.749617e-10, -2.742822e-10, -3.027227e-10, 
    -3.215591e-10, -4.916761e-10, -2.973536e-10, -2.446458e-10, 
    -2.828466e-10, -1.743664e-10, -2.818864e-10, -2.327283e-10, 
    -3.910147e-10, -3.419322e-10, -3.502926e-10, -3.865156e-10, 
    -3.319456e-10, -2.331425e-10, -4.738118e-10, -5.505583e-10, 
    -4.887333e-10, -4.353266e-10, -2.78589e-10, -3.018966e-10, -3.132332e-10, 
    -4.793209e-10, -4.673257e-10, -1.416687e-10, -4.392371e-10, 
    -3.837849e-10, -3.266865e-10, -1.764112e-10, -2.399062e-10, -2.40078e-10, 
    -3.205592e-10, -1.843672e-10, -2.875389e-10, -3.33184e-10, -4.197972e-10, 
    -2.613585e-10, -6.197909e-10, -2.788363e-10, -3.436621e-10, 
    -2.585336e-10, -3.358606e-10, -1.584903e-10, -2.072678e-10, 
    -3.524834e-10, -3.6909e-10, -3.739166e-10, -2.538238e-10, -4.770512e-10, 
    -3.724062e-10, -3.372659e-10, -2.087561e-10, -4.238355e-10, 
    -2.699774e-10, -3.461161e-10, -2.383662e-10, -3.544845e-10, -3.90739e-10, 
    -1.182698e-10, -1.437237e-10, -4.065989e-10, -3.367681e-10, 
    -2.108849e-10, -3.985659e-10, -3.586267e-10, -3.788161e-10, 
    -2.993126e-10, -5.636706e-10, -2.860789e-10, -2.940015e-10, 
    -4.980413e-10, -3.413944e-10, -3.916496e-10, -2.347496e-10, -3.58393e-10, 
    -1.874457e-10, -4.518163e-10, -2.956086e-10, -2.348246e-10, 
    -3.867575e-10, -3.404413e-10, -2.664231e-10, -2.305068e-10, 
    -2.472656e-10, -2.240705e-10, -2.677551e-10, -5.150683e-10, 
    -4.918954e-10, -4.689629e-10, -3.127162e-10, -4.527615e-10, 
    -4.647943e-10, -3.918421e-10, -3.780363e-10, -4.790849e-10, 
    -4.961278e-10, -2.595171e-10, -4.861958e-10, -2.217947e-10, 
    -3.452292e-10, -4.466309e-10, -3.281292e-10, -5.671141e-10, -4.13655e-10, 
    -1.894786e-10, -1.559887e-10, -2.978087e-10, -1.093896e-10, 
    -1.454277e-10, -1.977709e-10, -2.879975e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  5.976154e-16, 5.914084e-16, 5.926169e-16, 5.875984e-16, 5.903843e-16, 
    5.870955e-16, 5.963591e-16, 5.911611e-16, 5.944813e-16, 5.970581e-16, 
    5.778206e-16, 5.873744e-16, 5.6785e-16, 5.739805e-16, 5.585494e-16, 
    5.688043e-16, 5.564756e-16, 5.588471e-16, 5.517041e-16, 5.53753e-16, 
    5.445877e-16, 5.507578e-16, 5.398229e-16, 5.460635e-16, 5.450879e-16, 
    5.509608e-16, 5.854565e-16, 5.790122e-16, 5.858374e-16, 5.8492e-16, 
    5.85332e-16, 5.903264e-16, 5.928376e-16, 5.980896e-16, 5.971375e-16, 
    5.932799e-16, 5.845074e-16, 5.874905e-16, 5.799657e-16, 5.80136e-16, 
    5.717246e-16, 5.755215e-16, 5.613294e-16, 5.653729e-16, 5.536675e-16, 
    5.566174e-16, 5.53806e-16, 5.54659e-16, 5.537949e-16, 5.581195e-16, 
    5.562677e-16, 5.600695e-16, 5.748107e-16, 5.704878e-16, 5.833485e-16, 
    5.91038e-16, 5.961312e-16, 5.997362e-16, 5.99227e-16, 5.982556e-16, 
    5.932573e-16, 5.885468e-16, 5.849489e-16, 5.825384e-16, 5.801605e-16, 
    5.729421e-16, 5.691114e-16, 5.605102e-16, 5.620661e-16, 5.594304e-16, 
    5.569107e-16, 5.52672e-16, 5.533704e-16, 5.515007e-16, 5.595007e-16, 
    5.541869e-16, 5.629516e-16, 5.60558e-16, 5.795097e-16, 5.866863e-16, 
    5.897254e-16, 5.923845e-16, 5.988353e-16, 5.943827e-16, 5.961391e-16, 
    5.919585e-16, 5.892969e-16, 5.906139e-16, 5.824724e-16, 5.856415e-16, 
    5.688842e-16, 5.761208e-16, 5.572047e-16, 5.61747e-16, 5.561147e-16, 
    5.589908e-16, 5.5406e-16, 5.584982e-16, 5.508047e-16, 5.491252e-16, 
    5.502729e-16, 5.45862e-16, 5.587439e-16, 5.538057e-16, 5.906506e-16, 
    5.904359e-16, 5.894355e-16, 5.938289e-16, 5.940977e-16, 5.981156e-16, 
    5.945412e-16, 5.930167e-16, 5.891428e-16, 5.868469e-16, 5.846622e-16, 
    5.798502e-16, 5.744613e-16, 5.669003e-16, 5.614528e-16, 5.577929e-16, 
    5.600381e-16, 5.58056e-16, 5.602715e-16, 5.613093e-16, 5.497544e-16, 
    5.562502e-16, 5.464969e-16, 5.47038e-16, 5.51456e-16, 5.46977e-16, 
    5.902851e-16, 5.915206e-16, 5.958028e-16, 5.924524e-16, 5.985527e-16, 
    5.9514e-16, 5.931746e-16, 5.855745e-16, 5.839016e-16, 5.823479e-16, 
    5.792766e-16, 5.753273e-16, 5.683782e-16, 5.623146e-16, 5.567641e-16, 
    5.571714e-16, 5.57028e-16, 5.557858e-16, 5.58861e-16, 5.552805e-16, 
    5.546787e-16, 5.562514e-16, 5.471104e-16, 5.49726e-16, 5.470495e-16, 
    5.48753e-16, 5.911191e-16, 5.890396e-16, 5.901635e-16, 5.880492e-16, 
    5.895387e-16, 5.829057e-16, 5.809126e-16, 5.715605e-16, 5.754049e-16, 
    5.69282e-16, 5.747843e-16, 5.738106e-16, 5.690804e-16, 5.744878e-16, 
    5.626487e-16, 5.7068e-16, 5.557375e-16, 5.637832e-16, 5.552322e-16, 
    5.567882e-16, 5.542117e-16, 5.51901e-16, 5.489912e-16, 5.436104e-16, 
    5.448578e-16, 5.403509e-16, 5.859355e-16, 5.832301e-16, 5.834692e-16, 
    5.806348e-16, 5.785358e-16, 5.739795e-16, 5.666471e-16, 5.69407e-16, 
    5.643381e-16, 5.633188e-16, 5.710189e-16, 5.662939e-16, 5.81418e-16, 
    5.789819e-16, 5.804332e-16, 5.857218e-16, 5.687703e-16, 5.774887e-16, 
    5.613625e-16, 5.661066e-16, 5.522305e-16, 5.591423e-16, 5.45544e-16, 
    5.397022e-16, 5.341932e-16, 5.277338e-16, 5.817528e-16, 5.835928e-16, 
    5.802977e-16, 5.757282e-16, 5.71479e-16, 5.658174e-16, 5.652377e-16, 
    5.641748e-16, 5.614198e-16, 5.591002e-16, 5.638379e-16, 5.585184e-16, 
    5.78415e-16, 5.680124e-16, 5.842873e-16, 5.794003e-16, 5.759981e-16, 
    5.77492e-16, 5.697224e-16, 5.67887e-16, 5.604112e-16, 5.642796e-16, 
    5.411448e-16, 5.514116e-16, 5.228054e-16, 5.308367e-16, 5.842351e-16, 
    5.817595e-16, 5.73118e-16, 5.772345e-16, 5.654393e-16, 5.625255e-16, 
    5.601543e-16, 5.571181e-16, 5.567906e-16, 5.549894e-16, 5.579401e-16, 
    5.551063e-16, 5.658054e-16, 5.610312e-16, 5.741086e-16, 5.709314e-16, 
    5.72395e-16, 5.739964e-16, 5.690477e-16, 5.637632e-16, 5.636513e-16, 
    5.619535e-16, 5.571598e-16, 5.653914e-16, 5.398139e-16, 5.556448e-16, 
    5.790563e-16, 5.742709e-16, 5.735878e-16, 5.754433e-16, 5.628178e-16, 
    5.674007e-16, 5.550335e-16, 5.583835e-16, 5.52892e-16, 5.556225e-16, 
    5.560239e-16, 5.595252e-16, 5.617017e-16, 5.671906e-16, 5.71648e-16, 
    5.751745e-16, 5.743551e-16, 5.704774e-16, 5.634398e-16, 5.567604e-16, 
    5.582252e-16, 5.533099e-16, 5.662967e-16, 5.608604e-16, 5.629629e-16, 
    5.574765e-16, 5.6948e-16, 5.592593e-16, 5.720859e-16, 5.709629e-16, 
    5.674916e-16, 5.604904e-16, 5.589399e-16, 5.572811e-16, 5.583051e-16, 
    5.63261e-16, 5.640723e-16, 5.675763e-16, 5.685422e-16, 5.712072e-16, 
    5.734123e-16, 5.713972e-16, 5.692806e-16, 5.632594e-16, 5.578173e-16, 
    5.51868e-16, 5.504099e-16, 5.434296e-16, 5.49112e-16, 5.397252e-16, 
    5.477059e-16, 5.338735e-16, 5.586671e-16, 5.479425e-16, 5.673339e-16, 
    5.652539e-16, 5.61485e-16, 5.528172e-16, 5.575024e-16, 5.520226e-16, 
    5.641041e-16, 5.70343e-16, 5.719575e-16, 5.7496e-16, 5.718887e-16, 
    5.721388e-16, 5.691938e-16, 5.7014e-16, 5.630592e-16, 5.668658e-16, 
    5.560337e-16, 5.520663e-16, 5.408232e-16, 5.33901e-16, 5.268342e-16, 
    5.237066e-16, 5.227539e-16, 5.223555e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGR =
  -396.5523, -397.5788, -397.3809, -398.2022, -397.7469, -398.2845, 
    -396.7592, -397.619, -397.0677, -396.6445, -399.7943, -398.239, 
    -401.4218, -400.42, -402.921, -401.2672, -403.2544, -402.874, -404.0204, 
    -403.6921, -405.1562, -404.1719, -405.9157, -404.9215, -405.0768, 
    -404.1393, -398.5527, -399.6006, -398.4904, -398.6399, -398.573, 
    -397.7561, -397.3438, -396.4749, -396.6314, -397.2719, -398.7072, 
    -398.2205, -399.4481, -399.4204, -400.7858, -400.1703, -402.4746, 
    -401.823, -403.7058, -403.2324, -403.6835, -403.5468, -403.6852, 
    -402.9909, -403.2884, -402.6775, -400.2854, -400.9957, -398.8965, 
    -397.6384, -396.7965, -396.2037, -396.2875, -396.4472, -397.2756, 
    -398.0477, -398.6358, -399.029, -399.4164, -400.5869, -401.2179, 
    -402.606, -402.3561, -402.7798, -403.1853, -403.8651, -403.7534, 
    -404.0526, -402.7691, -403.622, -402.2137, -402.5989, -399.5195, 
    -398.3519, -397.8535, -397.4189, -396.3519, -397.0835, -396.7951, 
    -397.4891, -397.925, -397.7095, -399.0397, -398.5226, -401.2546, 
    -400.0725, -403.138, -402.4074, -403.3132, -402.8512, -403.6425, 
    -402.9304, -404.1642, -404.4325, -404.2491, -404.9543, -402.8908, 
    -403.6833, -397.7034, -397.7385, -397.9024, -397.1818, -397.1304, 
    -396.4705, -397.0579, -397.3152, -397.9504, -398.3256, -398.6824, 
    -399.4666, -400.3417, -401.5757, -402.4548, -403.0437, -402.6828, 
    -403.0014, -402.6451, -402.4782, -404.3318, -403.291, -404.8528, 
    -404.7665, -404.0597, -404.7763, -397.7632, -397.561, -396.8506, 
    -397.4082, -396.3986, -396.9593, -397.2889, -398.5329, -398.8067, 
    -399.0598, -399.5601, -400.2018, -401.337, -402.3157, -403.209, 
    -403.1436, -403.1666, -403.3659, -402.8719, -403.447, -403.5432, 
    -403.2912, -404.755, -404.3369, -404.7647, -404.4926, -397.6268, 
    -397.9671, -397.7832, -398.1289, -397.8852, -398.9682, -399.2928, 
    -400.8116, -400.189, -401.1907, -400.2899, -400.4476, -401.2221, 
    -400.3382, -402.2613, -400.9637, -403.3736, -402.0778, -403.4547, 
    -403.2051, -403.6186, -403.9886, -404.4544, -405.3128, -405.1142, 
    -405.8322, -398.4746, -398.9157, -398.8773, -399.3391, -399.6804, 
    -400.4206, -401.6169, -401.1711, -401.99, -402.1542, -400.9103, 
    -401.6737, -399.2112, -399.6071, -399.3717, -398.5092, -401.2733, 
    -399.85, -402.4692, -401.7044, -403.9358, -402.826, -405.0047, -405.9341, 
    -406.8104, -407.8314, -399.1568, -398.8571, -399.3941, -400.136, 
    -400.8355, -401.7509, -401.8448, -402.0161, -402.4604, -402.8335, 
    -402.0699, -402.9271, -399.6981, -401.3961, -398.7434, -399.5389, 
    -400.0924, -399.8501, -401.1203, -401.417, -402.6221, -401.9995, 
    -405.7044, -404.0662, -408.6099, -407.3411, -398.7523, -399.156, 
    -400.5597, -399.892, -401.8123, -402.282, -402.6641, -403.1517, 
    -403.2047, -403.4936, -403.0201, -403.475, -401.7529, -402.5227, 
    -400.3998, -400.9242, -400.6776, -400.418, -401.2293, -402.0818, 
    -402.1007, -402.3738, -403.1421, -401.82, -405.9144, -403.3858, 
    -399.5961, -400.3723, -400.4839, -400.1832, -402.2349, -401.4953, 
    -403.4866, -402.9488, -403.8301, -403.3922, -403.3277, -402.7652, 
    -402.4147, -401.5291, -400.7982, -400.2269, -400.3598, -400.9975, 
    -402.1341, -403.2091, -402.9736, -403.7632, -401.6738, -402.5498, 
    -402.2111, -403.0944, -401.1591, -402.8051, -400.7277, -400.9194, 
    -401.4806, -402.6088, -402.8593, -403.1255, -402.9614, -402.1631, 
    -402.0325, -401.4672, -401.3107, -400.8799, -400.5127, -400.8489, 
    -401.1911, -402.1637, -403.0393, -403.9938, -404.2275, -405.3401, 
    -404.4335, -405.9284, -404.6562, -406.8586, -402.9015, -404.6201, 
    -401.5064, -401.8423, -402.4489, -403.8409, -403.0902, -403.9684, 
    -402.0275, -401.0188, -400.7484, -400.2615, -400.7596, -400.7191, 
    -401.2058, -401.0527, -402.196, -401.582, -403.3259, -403.9616, 
    -405.7567, -406.8557, -407.9748, -408.4682, -408.6184, -408.6812 ;

 FGR12 =
  -51.97826, -52.04658, -52.03333, -52.08843, -52.0579, -52.09396, -51.99214, 
    -52.04925, -52.01281, -51.98446, -52.19544, -52.09092, -52.30472, 
    -52.23777, -52.40617, -52.29428, -52.4288, -52.40306, -52.48083, 
    -52.45855, -52.55795, -52.49114, -52.6097, -52.54205, -52.55257, 
    -52.48892, -52.11203, -52.18239, -52.10783, -52.11787, -52.11337, 
    -52.05849, -52.03077, -51.9731, -51.98358, -52.02599, -52.12238, 
    -52.08971, -52.17229, -52.17043, -52.26245, -52.22095, -52.376, 
    -52.33192, -52.45947, -52.42736, -52.45795, -52.44869, -52.45807, 
    -52.41098, -52.43114, -52.38975, -52.22869, -52.27597, -52.13512, 
    -52.05053, -51.99462, -51.95494, -51.96054, -51.97121, -52.02624, 
    -52.07809, -52.11763, -52.14407, -52.17017, -52.24894, -52.29097, 
    -52.38486, -52.368, -52.39665, -52.42417, -52.47027, -52.4627, -52.483, 
    -52.39597, -52.45376, -52.35836, -52.38442, -52.17692, -52.09854, 
    -52.06497, -52.03586, -51.96486, -52.01384, -51.99452, -52.04059, 
    -52.06985, -52.0554, -52.14479, -52.11001, -52.29343, -52.21433, 
    -52.42094, -52.37146, -52.43283, -52.40153, -52.45516, -52.40689, 
    -52.49059, -52.5088, -52.49635, -52.54428, -52.40421, -52.45792, 
    -52.05498, -52.05733, -52.06833, -52.01995, -52.01699, -51.9728, 
    -52.01215, -52.0289, -52.07157, -52.09676, -52.12075, -52.17351, 
    -52.23248, -52.31515, -52.37467, -52.41457, -52.39012, -52.4117, 
    -52.38757, -52.37627, -52.50195, -52.43132, -52.5374, -52.53154, 
    -52.48348, -52.53218, -52.05899, -52.04543, -51.99826, -52.03516, 
    -51.96799, -52.00553, -52.02713, -52.11065, -52.12912, -52.14613, 
    -52.17983, -52.22306, -52.29904, -52.36522, -52.42578, -52.42134, 
    -52.4229, -52.43641, -52.40293, -52.4419, -52.44842, -52.43135, 
    -52.53074, -52.50233, -52.53141, -52.51292, -52.04985, -52.07268, 
    -52.06034, -52.08354, -52.06717, -52.13992, -52.16178, -52.26414, 
    -52.2222, -52.28913, -52.22901, -52.23963, -52.29119, -52.23228, 
    -52.3615, -52.27378, -52.43692, -52.34907, -52.44243, -52.42552, 
    -52.45356, -52.47866, -52.51032, -52.56866, -52.55517, -52.60405, 
    -52.10679, -52.13641, -52.13387, -52.16493, -52.18792, -52.23782, 
    -52.31796, -52.28786, -52.34321, -52.35431, -52.27026, -52.32179, 
    -52.15631, -52.18293, -52.16712, -52.1091, -52.2947, -52.19932, 
    -52.37563, -52.32389, -52.47507, -52.39978, -52.54772, -52.61092, 
    -52.67078, -52.74046, -52.15266, -52.13252, -52.16866, -52.21858, 
    -52.26519, -52.32702, -52.3334, -52.34497, -52.37505, -52.40033, 
    -52.34858, -52.40666, -52.18901, -52.30301, -52.12486, -52.17833, 
    -52.21567, -52.19935, -52.28444, -52.30447, -52.38597, -52.34386, 
    -52.59526, -52.48389, -52.79377, -52.70697, -52.12547, -52.15262, 
    -52.24718, -52.20218, -52.33119, -52.36296, -52.38885, -52.42187, 
    -52.42548, -52.44506, -52.41297, -52.44381, -52.32717, -52.37926, 
    -52.23644, -52.27117, -52.25517, -52.23766, -52.29181, -52.34937, 
    -52.35071, -52.36916, -52.42104, -52.33174, -52.60946, -52.43763, 
    -52.18226, -52.2345, -52.24209, -52.22182, -52.35977, -52.30976, 
    -52.44459, -52.40814, -52.4679, -52.4382, -52.43381, -52.3957, -52.37194, 
    -52.31203, -52.26329, -52.22478, -52.23374, -52.27611, -52.35293, 
    -52.42575, -52.40979, -52.46336, -52.32185, -52.38108, -52.35816, 
    -52.418, -52.28705, -52.39822, -52.25856, -52.27087, -52.30877, 
    -52.38503, -52.40208, -52.42009, -52.40899, -52.3549, -52.34608, 
    -52.30787, -52.29726, -52.26821, -52.24406, -52.2661, -52.28919, 
    -52.35495, -52.41426, -52.47899, -52.49491, -52.57043, -52.50882, 
    -52.61041, -52.52385, -52.67391, -52.40485, -52.52145, -52.31053, 
    -52.33323, -52.37423, -52.46856, -52.41772, -52.47724, -52.34574, 
    -52.27753, -52.25995, -52.22711, -52.26071, -52.25798, -52.29021, 
    -52.27987, -52.35714, -52.31563, -52.43369, -52.4768, -52.5989, 
    -52.67381, -52.75033, -52.78411, -52.79439, -52.7987 ;

 FGR_R =
  -396.5523, -397.5788, -397.3809, -398.2022, -397.7469, -398.2845, 
    -396.7592, -397.619, -397.0677, -396.6445, -399.7943, -398.239, 
    -401.4218, -400.42, -402.921, -401.2672, -403.2544, -402.874, -404.0204, 
    -403.6921, -405.1562, -404.1719, -405.9157, -404.9215, -405.0768, 
    -404.1393, -398.5527, -399.6006, -398.4904, -398.6399, -398.573, 
    -397.7561, -397.3438, -396.4749, -396.6314, -397.2719, -398.7072, 
    -398.2205, -399.4481, -399.4204, -400.7858, -400.1703, -402.4746, 
    -401.823, -403.7058, -403.2324, -403.6835, -403.5468, -403.6852, 
    -402.9909, -403.2884, -402.6775, -400.2854, -400.9957, -398.8965, 
    -397.6384, -396.7965, -396.2037, -396.2875, -396.4472, -397.2756, 
    -398.0477, -398.6358, -399.029, -399.4164, -400.5869, -401.2179, 
    -402.606, -402.3561, -402.7798, -403.1853, -403.8651, -403.7534, 
    -404.0526, -402.7691, -403.622, -402.2137, -402.5989, -399.5195, 
    -398.3519, -397.8535, -397.4189, -396.3519, -397.0835, -396.7951, 
    -397.4891, -397.925, -397.7095, -399.0397, -398.5226, -401.2546, 
    -400.0725, -403.138, -402.4074, -403.3132, -402.8512, -403.6425, 
    -402.9304, -404.1642, -404.4325, -404.2491, -404.9543, -402.8908, 
    -403.6833, -397.7034, -397.7385, -397.9024, -397.1818, -397.1304, 
    -396.4705, -397.0579, -397.3152, -397.9504, -398.3256, -398.6824, 
    -399.4666, -400.3417, -401.5757, -402.4548, -403.0437, -402.6828, 
    -403.0014, -402.6451, -402.4782, -404.3318, -403.291, -404.8528, 
    -404.7665, -404.0597, -404.7763, -397.7632, -397.561, -396.8506, 
    -397.4082, -396.3986, -396.9593, -397.2889, -398.5329, -398.8067, 
    -399.0598, -399.5601, -400.2018, -401.337, -402.3157, -403.209, 
    -403.1436, -403.1666, -403.3659, -402.8719, -403.447, -403.5432, 
    -403.2912, -404.755, -404.3369, -404.7647, -404.4926, -397.6268, 
    -397.9671, -397.7832, -398.1289, -397.8852, -398.9682, -399.2928, 
    -400.8116, -400.189, -401.1907, -400.2899, -400.4476, -401.2221, 
    -400.3382, -402.2613, -400.9637, -403.3736, -402.0778, -403.4547, 
    -403.2051, -403.6186, -403.9886, -404.4544, -405.3128, -405.1142, 
    -405.8322, -398.4746, -398.9157, -398.8773, -399.3391, -399.6804, 
    -400.4206, -401.6169, -401.1711, -401.99, -402.1542, -400.9103, 
    -401.6737, -399.2112, -399.6071, -399.3717, -398.5092, -401.2733, 
    -399.85, -402.4692, -401.7044, -403.9358, -402.826, -405.0047, -405.9341, 
    -406.8104, -407.8314, -399.1568, -398.8571, -399.3941, -400.136, 
    -400.8355, -401.7509, -401.8448, -402.0161, -402.4604, -402.8335, 
    -402.0699, -402.9271, -399.6981, -401.3961, -398.7434, -399.5389, 
    -400.0924, -399.8501, -401.1203, -401.417, -402.6221, -401.9995, 
    -405.7044, -404.0662, -408.6099, -407.3411, -398.7523, -399.156, 
    -400.5597, -399.892, -401.8123, -402.282, -402.6641, -403.1517, 
    -403.2047, -403.4936, -403.0201, -403.475, -401.7529, -402.5227, 
    -400.3998, -400.9242, -400.6776, -400.418, -401.2293, -402.0818, 
    -402.1007, -402.3738, -403.1421, -401.82, -405.9144, -403.3858, 
    -399.5961, -400.3723, -400.4839, -400.1832, -402.2349, -401.4953, 
    -403.4866, -402.9488, -403.8301, -403.3922, -403.3277, -402.7652, 
    -402.4147, -401.5291, -400.7982, -400.2269, -400.3598, -400.9975, 
    -402.1341, -403.2091, -402.9736, -403.7632, -401.6738, -402.5498, 
    -402.2111, -403.0944, -401.1591, -402.8051, -400.7277, -400.9194, 
    -401.4806, -402.6088, -402.8593, -403.1255, -402.9614, -402.1631, 
    -402.0325, -401.4672, -401.3107, -400.8799, -400.5127, -400.8489, 
    -401.1911, -402.1637, -403.0393, -403.9938, -404.2275, -405.3401, 
    -404.4335, -405.9284, -404.6562, -406.8586, -402.9015, -404.6201, 
    -401.5064, -401.8423, -402.4489, -403.8409, -403.0902, -403.9684, 
    -402.0275, -401.0188, -400.7484, -400.2615, -400.7596, -400.7191, 
    -401.2058, -401.0527, -402.196, -401.582, -403.3259, -403.9616, 
    -405.7567, -406.8557, -407.9748, -408.4682, -408.6184, -408.6812 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  48.64191, 48.7161, 48.70165, 48.76162, 48.72838, 48.76763, 48.65702, 
    48.71903, 48.67955, 48.64864, 48.87788, 48.76431, 48.99442, 48.9236, 
    49.10389, 48.98312, 49.12825, 49.10047, 49.18419, 49.16022, 49.26711, 
    49.19526, 49.32259, 49.24999, 49.26133, 49.19287, 48.78722, 48.86372, 
    48.78268, 48.79359, 48.78871, 48.72905, 48.69893, 48.63626, 48.64769, 
    48.69368, 48.7985, 48.76297, 48.85262, 48.8506, 48.95031, 48.90536, 
    49.0713, 49.02373, 49.16122, 49.12664, 49.15958, 49.1496, 49.15971, 
    49.10901, 49.13073, 49.08612, 48.91377, 48.96332, 48.81233, 48.72044, 
    48.65974, 48.61646, 48.62257, 48.63423, 48.69395, 48.75035, 48.7933, 
    48.82201, 48.85031, 48.93577, 48.97953, 49.08089, 49.06266, 49.09359, 
    49.12321, 49.17285, 49.16469, 49.18654, 49.09281, 49.15509, 49.05226, 
    49.08038, 48.8578, 48.77256, 48.73615, 48.70442, 48.62728, 48.6807, 
    48.65964, 48.70956, 48.74139, 48.72565, 48.8228, 48.78503, 48.98222, 
    48.89822, 49.11975, 49.06641, 49.13255, 49.09881, 49.15659, 49.10459, 
    49.19469, 49.21428, 49.20089, 49.25238, 49.1017, 49.15956, 48.7252, 
    48.72777, 48.73974, 48.68711, 48.68412, 48.63593, 48.67883, 48.69685, 
    48.74324, 48.77065, 48.7967, 48.85397, 48.91788, 49.00566, 49.06986, 
    49.11287, 49.08651, 49.10978, 49.08376, 49.07157, 49.20692, 49.13092, 
    49.24498, 49.23868, 49.18705, 49.23939, 48.72957, 48.71481, 48.66369, 
    48.70364, 48.63069, 48.67163, 48.69493, 48.78577, 48.80577, 48.82426, 
    48.8608, 48.90766, 48.98824, 49.0597, 49.12494, 49.12016, 49.12184, 
    49.13639, 49.10032, 49.14231, 49.14934, 49.13094, 49.23783, 49.20731, 
    49.23854, 49.21867, 48.71961, 48.74446, 48.73103, 48.75628, 48.73848, 
    48.81756, 48.84127, 48.95219, 48.90673, 48.97755, 48.9141, 48.92561, 
    48.97983, 48.91763, 49.05572, 48.96097, 49.13696, 49.04231, 49.14288, 
    49.12466, 49.15485, 49.18187, 49.21588, 49.27856, 49.26406, 49.31649, 
    48.78152, 48.81373, 48.81093, 48.84465, 48.86958, 48.92364, 49.00868, 
    48.97613, 49.03592, 49.04791, 48.95709, 49.01283, 48.83531, 48.86422, 
    48.84703, 48.78405, 48.98358, 48.88196, 49.07092, 49.01506, 49.17801, 
    49.09696, 49.25607, 49.32393, 49.38794, 49.46249, 48.83134, 48.80946, 
    48.84867, 48.90285, 48.95162, 49.01846, 49.02532, 49.03783, 49.07027, 
    49.09752, 49.04175, 49.10435, 48.87085, 48.99255, 48.80116, 48.85924, 
    48.89967, 48.88197, 48.97242, 48.99408, 49.08207, 49.03661, 49.30715, 
    49.18752, 49.51936, 49.42669, 48.80181, 48.83129, 48.9338, 48.88504, 
    49.02295, 49.05724, 49.08515, 49.12075, 49.12462, 49.14571, 49.11114, 
    49.14436, 49.01861, 49.07483, 48.92213, 48.9581, 48.94241, 48.92345, 
    48.98038, 49.04262, 49.04401, 49.06395, 49.12001, 49.02351, 49.32246, 
    49.13781, 48.86343, 48.9201, 48.92827, 48.9063, 49.0538, 48.9998, 
    49.14521, 49.10594, 49.17029, 49.13831, 49.1336, 49.09253, 49.06694, 
    49.00227, 48.95121, 48.9095, 48.9192, 48.96345, 49.04644, 49.12494, 
    49.10774, 49.1654, 49.01284, 49.0768, 49.05206, 49.11657, 48.97525, 
    49.09541, 48.94608, 48.95775, 48.99873, 49.08109, 49.0994, 49.11884, 
    49.10686, 49.04855, 49.03903, 48.99775, 48.98632, 48.95487, 48.93037, 
    48.95261, 48.97758, 49.0486, 49.11254, 49.18224, 49.19931, 49.28054, 
    49.21434, 49.32348, 49.23057, 49.39143, 49.10246, 49.22796, 49.00061, 
    49.02514, 49.06942, 49.17107, 49.11626, 49.18038, 49.03866, 48.965, 
    48.94759, 48.91203, 48.9484, 48.94545, 48.97866, 48.96749, 49.05096, 
    49.00613, 49.13347, 49.17989, 49.31098, 49.39124, 49.47298, 49.50901, 
    49.51999, 49.52457 ;

 FIRA_R =
  48.64191, 48.7161, 48.70165, 48.76162, 48.72838, 48.76763, 48.65702, 
    48.71903, 48.67955, 48.64864, 48.87788, 48.76431, 48.99442, 48.9236, 
    49.10389, 48.98312, 49.12825, 49.10047, 49.18419, 49.16022, 49.26711, 
    49.19526, 49.32259, 49.24999, 49.26133, 49.19287, 48.78722, 48.86372, 
    48.78268, 48.79359, 48.78871, 48.72905, 48.69893, 48.63626, 48.64769, 
    48.69368, 48.7985, 48.76297, 48.85262, 48.8506, 48.95031, 48.90536, 
    49.0713, 49.02373, 49.16122, 49.12664, 49.15958, 49.1496, 49.15971, 
    49.10901, 49.13073, 49.08612, 48.91377, 48.96332, 48.81233, 48.72044, 
    48.65974, 48.61646, 48.62257, 48.63423, 48.69395, 48.75035, 48.7933, 
    48.82201, 48.85031, 48.93577, 48.97953, 49.08089, 49.06266, 49.09359, 
    49.12321, 49.17285, 49.16469, 49.18654, 49.09281, 49.15509, 49.05226, 
    49.08038, 48.8578, 48.77256, 48.73615, 48.70442, 48.62728, 48.6807, 
    48.65964, 48.70956, 48.74139, 48.72565, 48.8228, 48.78503, 48.98222, 
    48.89822, 49.11975, 49.06641, 49.13255, 49.09881, 49.15659, 49.10459, 
    49.19469, 49.21428, 49.20089, 49.25238, 49.1017, 49.15956, 48.7252, 
    48.72777, 48.73974, 48.68711, 48.68412, 48.63593, 48.67883, 48.69685, 
    48.74324, 48.77065, 48.7967, 48.85397, 48.91788, 49.00566, 49.06986, 
    49.11287, 49.08651, 49.10978, 49.08376, 49.07157, 49.20692, 49.13092, 
    49.24498, 49.23868, 49.18705, 49.23939, 48.72957, 48.71481, 48.66369, 
    48.70364, 48.63069, 48.67163, 48.69493, 48.78577, 48.80577, 48.82426, 
    48.8608, 48.90766, 48.98824, 49.0597, 49.12494, 49.12016, 49.12184, 
    49.13639, 49.10032, 49.14231, 49.14934, 49.13094, 49.23783, 49.20731, 
    49.23854, 49.21867, 48.71961, 48.74446, 48.73103, 48.75628, 48.73848, 
    48.81756, 48.84127, 48.95219, 48.90673, 48.97755, 48.9141, 48.92561, 
    48.97983, 48.91763, 49.05572, 48.96097, 49.13696, 49.04231, 49.14288, 
    49.12466, 49.15485, 49.18187, 49.21588, 49.27856, 49.26406, 49.31649, 
    48.78152, 48.81373, 48.81093, 48.84465, 48.86958, 48.92364, 49.00868, 
    48.97613, 49.03592, 49.04791, 48.95709, 49.01283, 48.83531, 48.86422, 
    48.84703, 48.78405, 48.98358, 48.88196, 49.07092, 49.01506, 49.17801, 
    49.09696, 49.25607, 49.32393, 49.38794, 49.46249, 48.83134, 48.80946, 
    48.84867, 48.90285, 48.95162, 49.01846, 49.02532, 49.03783, 49.07027, 
    49.09752, 49.04175, 49.10435, 48.87085, 48.99255, 48.80116, 48.85924, 
    48.89967, 48.88197, 48.97242, 48.99408, 49.08207, 49.03661, 49.30715, 
    49.18752, 49.51936, 49.42669, 48.80181, 48.83129, 48.9338, 48.88504, 
    49.02295, 49.05724, 49.08515, 49.12075, 49.12462, 49.14571, 49.11114, 
    49.14436, 49.01861, 49.07483, 48.92213, 48.9581, 48.94241, 48.92345, 
    48.98038, 49.04262, 49.04401, 49.06395, 49.12001, 49.02351, 49.32246, 
    49.13781, 48.86343, 48.9201, 48.92827, 48.9063, 49.0538, 48.9998, 
    49.14521, 49.10594, 49.17029, 49.13831, 49.1336, 49.09253, 49.06694, 
    49.00227, 48.95121, 48.9095, 48.9192, 48.96345, 49.04644, 49.12494, 
    49.10774, 49.1654, 49.01284, 49.0768, 49.05206, 49.11657, 48.97525, 
    49.09541, 48.94608, 48.95775, 48.99873, 49.08109, 49.0994, 49.11884, 
    49.10686, 49.04855, 49.03903, 48.99775, 48.98632, 48.95487, 48.93037, 
    48.95261, 48.97758, 49.0486, 49.11254, 49.18224, 49.19931, 49.28054, 
    49.21434, 49.32348, 49.23057, 49.39143, 49.10246, 49.22796, 49.00061, 
    49.02514, 49.06942, 49.17107, 49.11626, 49.18038, 49.03866, 48.965, 
    48.94759, 48.91203, 48.9484, 48.94545, 48.97866, 48.96749, 49.05096, 
    49.00613, 49.13347, 49.17989, 49.31098, 49.39124, 49.47298, 49.50901, 
    49.51999, 49.52457 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  262.988, 263.0623, 263.0478, 263.1078, 263.0745, 263.1138, 263.0032, 
    263.0652, 263.0257, 262.9948, 263.224, 263.1104, 263.3406, 263.2697, 
    263.45, 263.3293, 263.4744, 263.4466, 263.5303, 263.5063, 263.6133, 
    263.5414, 263.6687, 263.5961, 263.6075, 263.539, 263.1334, 263.2099, 
    263.1288, 263.1397, 263.1349, 263.0752, 263.0451, 262.9824, 262.9938, 
    263.0398, 263.1447, 263.1091, 263.1988, 263.1967, 263.2964, 263.2515, 
    263.4174, 263.3699, 263.5074, 263.4728, 263.5057, 263.4958, 263.5059, 
    263.4551, 263.4769, 263.4323, 263.2599, 263.3094, 263.1585, 263.0666, 
    263.0059, 262.9626, 262.9687, 262.9804, 263.0401, 263.0965, 263.1394, 
    263.1682, 263.1964, 263.2819, 263.3257, 263.427, 263.4088, 263.4397, 
    263.4694, 263.519, 263.5108, 263.5327, 263.439, 263.5013, 263.3984, 
    263.4265, 263.2039, 263.1187, 263.0823, 263.0506, 262.9734, 263.0269, 
    263.0058, 263.0557, 263.0875, 263.0718, 263.1689, 263.1312, 263.3284, 
    263.2444, 263.4659, 263.4125, 263.4787, 263.4449, 263.5027, 263.4507, 
    263.5408, 263.5604, 263.547, 263.5985, 263.4478, 263.5057, 263.0714, 
    263.0739, 263.0859, 263.0333, 263.0303, 262.9821, 263.025, 263.043, 
    263.0894, 263.1168, 263.1429, 263.2001, 263.264, 263.3518, 263.416, 
    263.459, 263.4326, 263.4559, 263.4299, 263.4177, 263.5531, 263.4771, 
    263.5911, 263.5848, 263.5332, 263.5855, 263.0757, 263.0609, 263.0098, 
    263.0498, 262.9768, 263.0178, 263.0411, 263.1319, 263.1519, 263.1704, 
    263.2069, 263.2538, 263.3344, 263.4059, 263.4711, 263.4663, 263.468, 
    263.4825, 263.4465, 263.4885, 263.4955, 263.4771, 263.584, 263.5534, 
    263.5847, 263.5648, 263.0658, 263.0906, 263.0772, 263.1024, 263.0846, 
    263.1637, 263.1874, 263.2983, 263.2529, 263.3237, 263.2603, 263.2718, 
    263.326, 263.2638, 263.4019, 263.3071, 263.4831, 263.3885, 263.489, 
    263.4708, 263.501, 263.528, 263.562, 263.6247, 263.6102, 263.6626, 
    263.1277, 263.1599, 263.1571, 263.1908, 263.2157, 263.2698, 263.3548, 
    263.3223, 263.3821, 263.394, 263.3032, 263.359, 263.1815, 263.2104, 
    263.1932, 263.1302, 263.3297, 263.2281, 263.4171, 263.3612, 263.5241, 
    263.4431, 263.6022, 263.6701, 263.7341, 263.8086, 263.1775, 263.1556, 
    263.1948, 263.249, 263.2978, 263.3646, 263.3715, 263.384, 263.4164, 
    263.4437, 263.3879, 263.4505, 263.217, 263.3387, 263.1473, 263.2054, 
    263.2458, 263.2281, 263.3186, 263.3402, 263.4282, 263.3828, 263.6533, 
    263.5337, 263.8655, 263.7728, 263.1479, 263.1774, 263.2799, 263.2312, 
    263.3691, 263.4034, 263.4313, 263.4669, 263.4708, 263.4919, 263.4573, 
    263.4905, 263.3647, 263.421, 263.2683, 263.3042, 263.2885, 263.2696, 
    263.3265, 263.3888, 263.3901, 263.4101, 263.4662, 263.3697, 263.6686, 
    263.4839, 263.2096, 263.2662, 263.2744, 263.2524, 263.3999, 263.3459, 
    263.4914, 263.4521, 263.5164, 263.4845, 263.4797, 263.4387, 263.4131, 
    263.3484, 263.2974, 263.2556, 263.2654, 263.3096, 263.3926, 263.4711, 
    263.4539, 263.5115, 263.359, 263.4229, 263.3982, 263.4627, 263.3214, 
    263.4416, 263.2922, 263.3039, 263.3449, 263.4272, 263.4456, 263.465, 
    263.453, 263.3947, 263.3852, 263.3439, 263.3325, 263.301, 263.2765, 
    263.2987, 263.3237, 263.3947, 263.4587, 263.5284, 263.5455, 263.6267, 
    263.5605, 263.6696, 263.5767, 263.7376, 263.4486, 263.5741, 263.3468, 
    263.3713, 263.4156, 263.5172, 263.4624, 263.5265, 263.3848, 263.3112, 
    263.2937, 263.2582, 263.2946, 263.2916, 263.3248, 263.3136, 263.3971, 
    263.3523, 263.4796, 263.526, 263.6571, 263.7374, 263.8191, 263.8552, 
    263.8661, 263.8707 ;

 FIRE_R =
  262.988, 263.0623, 263.0478, 263.1078, 263.0745, 263.1138, 263.0032, 
    263.0652, 263.0257, 262.9948, 263.224, 263.1104, 263.3406, 263.2697, 
    263.45, 263.3293, 263.4744, 263.4466, 263.5303, 263.5063, 263.6133, 
    263.5414, 263.6687, 263.5961, 263.6075, 263.539, 263.1334, 263.2099, 
    263.1288, 263.1397, 263.1349, 263.0752, 263.0451, 262.9824, 262.9938, 
    263.0398, 263.1447, 263.1091, 263.1988, 263.1967, 263.2964, 263.2515, 
    263.4174, 263.3699, 263.5074, 263.4728, 263.5057, 263.4958, 263.5059, 
    263.4551, 263.4769, 263.4323, 263.2599, 263.3094, 263.1585, 263.0666, 
    263.0059, 262.9626, 262.9687, 262.9804, 263.0401, 263.0965, 263.1394, 
    263.1682, 263.1964, 263.2819, 263.3257, 263.427, 263.4088, 263.4397, 
    263.4694, 263.519, 263.5108, 263.5327, 263.439, 263.5013, 263.3984, 
    263.4265, 263.2039, 263.1187, 263.0823, 263.0506, 262.9734, 263.0269, 
    263.0058, 263.0557, 263.0875, 263.0718, 263.1689, 263.1312, 263.3284, 
    263.2444, 263.4659, 263.4125, 263.4787, 263.4449, 263.5027, 263.4507, 
    263.5408, 263.5604, 263.547, 263.5985, 263.4478, 263.5057, 263.0714, 
    263.0739, 263.0859, 263.0333, 263.0303, 262.9821, 263.025, 263.043, 
    263.0894, 263.1168, 263.1429, 263.2001, 263.264, 263.3518, 263.416, 
    263.459, 263.4326, 263.4559, 263.4299, 263.4177, 263.5531, 263.4771, 
    263.5911, 263.5848, 263.5332, 263.5855, 263.0757, 263.0609, 263.0098, 
    263.0498, 262.9768, 263.0178, 263.0411, 263.1319, 263.1519, 263.1704, 
    263.2069, 263.2538, 263.3344, 263.4059, 263.4711, 263.4663, 263.468, 
    263.4825, 263.4465, 263.4885, 263.4955, 263.4771, 263.584, 263.5534, 
    263.5847, 263.5648, 263.0658, 263.0906, 263.0772, 263.1024, 263.0846, 
    263.1637, 263.1874, 263.2983, 263.2529, 263.3237, 263.2603, 263.2718, 
    263.326, 263.2638, 263.4019, 263.3071, 263.4831, 263.3885, 263.489, 
    263.4708, 263.501, 263.528, 263.562, 263.6247, 263.6102, 263.6626, 
    263.1277, 263.1599, 263.1571, 263.1908, 263.2157, 263.2698, 263.3548, 
    263.3223, 263.3821, 263.394, 263.3032, 263.359, 263.1815, 263.2104, 
    263.1932, 263.1302, 263.3297, 263.2281, 263.4171, 263.3612, 263.5241, 
    263.4431, 263.6022, 263.6701, 263.7341, 263.8086, 263.1775, 263.1556, 
    263.1948, 263.249, 263.2978, 263.3646, 263.3715, 263.384, 263.4164, 
    263.4437, 263.3879, 263.4505, 263.217, 263.3387, 263.1473, 263.2054, 
    263.2458, 263.2281, 263.3186, 263.3402, 263.4282, 263.3828, 263.6533, 
    263.5337, 263.8655, 263.7728, 263.1479, 263.1774, 263.2799, 263.2312, 
    263.3691, 263.4034, 263.4313, 263.4669, 263.4708, 263.4919, 263.4573, 
    263.4905, 263.3647, 263.421, 263.2683, 263.3042, 263.2885, 263.2696, 
    263.3265, 263.3888, 263.3901, 263.4101, 263.4662, 263.3697, 263.6686, 
    263.4839, 263.2096, 263.2662, 263.2744, 263.2524, 263.3999, 263.3459, 
    263.4914, 263.4521, 263.5164, 263.4845, 263.4797, 263.4387, 263.4131, 
    263.3484, 263.2974, 263.2556, 263.2654, 263.3096, 263.3926, 263.4711, 
    263.4539, 263.5115, 263.359, 263.4229, 263.3982, 263.4627, 263.3214, 
    263.4416, 263.2922, 263.3039, 263.3449, 263.4272, 263.4456, 263.465, 
    263.453, 263.3947, 263.3852, 263.3439, 263.3325, 263.301, 263.2765, 
    263.2987, 263.3237, 263.3947, 263.4587, 263.5284, 263.5455, 263.6267, 
    263.5605, 263.6696, 263.5767, 263.7376, 263.4486, 263.5741, 263.3468, 
    263.3713, 263.4156, 263.5172, 263.4624, 263.5265, 263.3848, 263.3112, 
    263.2937, 263.2582, 263.2946, 263.2916, 263.3248, 263.3136, 263.3971, 
    263.3523, 263.4796, 263.526, 263.6571, 263.7374, 263.8191, 263.8552, 
    263.8661, 263.8707 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  347.9627, 348.915, 348.7315, 349.4929, 349.0708, 349.5691, 348.1545, 
    348.9522, 348.4404, 348.0481, 350.9688, 349.5269, 352.4797, 351.5487, 
    353.8694, 352.3363, 354.1785, 353.8258, 354.8885, 354.5842, 355.9413, 
    355.029, 356.6454, 355.7238, 355.8678, 354.9987, 349.8177, 350.7891, 
    349.76, 349.8986, 349.8366, 349.0793, 348.6972, 347.8909, 348.036, 
    348.6305, 349.961, 349.5098, 350.6478, 350.6221, 351.8878, 351.3172, 
    353.4556, 352.8515, 354.5969, 354.1581, 354.5762, 354.4495, 354.5778, 
    353.9342, 354.21, 353.6437, 351.424, 352.0847, 350.1364, 348.9702, 
    348.1891, 347.6396, 347.7173, 347.8652, 348.6339, 349.3497, 349.8948, 
    350.2593, 350.6184, 351.7034, 352.2906, 353.5774, 353.3458, 353.7385, 
    354.1144, 354.7446, 354.641, 354.9184, 353.7285, 354.5192, 353.2137, 
    353.5708, 350.714, 349.6317, 349.1696, 348.7667, 347.7769, 348.4551, 
    348.1878, 348.8318, 349.2359, 349.0362, 350.2693, 349.7899, 352.3247, 
    351.2266, 354.0706, 353.3933, 354.2329, 353.8047, 354.5382, 353.8781, 
    355.0218, 355.2705, 355.1005, 355.7542, 353.8414, 354.576, 349.0305, 
    349.063, 349.215, 348.5469, 348.4986, 347.8868, 348.4313, 348.6707, 
    349.2595, 349.6073, 349.938, 350.6649, 351.4761, 352.6223, 353.4372, 
    353.9831, 353.6486, 353.9439, 353.6136, 353.4589, 355.1772, 354.2124, 
    355.6602, 355.5802, 354.9249, 355.5892, 349.0859, 348.8985, 348.2392, 
    348.7568, 347.8202, 348.34, 348.6463, 349.7994, 350.0532, 350.2878, 
    350.7516, 351.3464, 352.401, 353.3083, 354.1364, 354.0757, 354.097, 
    354.2818, 353.8239, 354.357, 354.4462, 354.2125, 355.5694, 355.1819, 
    355.5785, 355.3262, 348.9595, 349.275, 349.1045, 349.425, 349.199, 
    350.2029, 350.5038, 351.9117, 351.3346, 352.2654, 351.4281, 351.5743, 
    352.2945, 351.4729, 353.2579, 352.0551, 354.2889, 353.0877, 354.3642, 
    354.1328, 354.5161, 354.859, 355.2908, 356.0865, 355.9024, 356.568, 
    349.7454, 350.1542, 350.1187, 350.5467, 350.8631, 351.5492, 352.6606, 
    352.2473, 353.0063, 353.1586, 352.0056, 352.7132, 350.4281, 350.7952, 
    350.5769, 349.7774, 352.342, 351.0203, 353.4506, 352.7416, 354.8101, 
    353.7813, 355.8009, 356.6625, 357.4747, 358.4212, 350.3778, 350.1, 
    350.5977, 351.2854, 351.9362, 352.7848, 352.8718, 353.0306, 353.4424, 
    353.7883, 353.0804, 353.875, 350.8795, 352.4558, 349.9946, 350.732, 
    351.2451, 351.0204, 352.2001, 352.4752, 353.5923, 353.0151, 356.4496, 
    354.9309, 359.1428, 357.9667, 350.0028, 350.377, 351.6782, 351.0593, 
    352.8416, 353.277, 353.6312, 354.0833, 354.1323, 354.4001, 353.9612, 
    354.3829, 352.7866, 353.5002, 351.53, 352.0184, 351.7875, 351.5468, 
    352.3012, 353.0915, 353.109, 353.3622, 354.0744, 352.8488, 356.6443, 
    354.3003, 350.7849, 351.5045, 351.608, 351.3292, 353.2333, 352.5478, 
    354.3937, 353.8951, 354.7121, 354.3062, 354.2464, 353.7249, 353.4001, 
    352.5791, 351.8992, 351.3697, 351.4929, 352.0864, 353.14, 354.1365, 
    353.9182, 354.65, 352.7133, 353.5253, 353.2113, 354.0301, 352.2362, 
    353.762, 351.8339, 352.0139, 352.5342, 353.58, 353.8122, 354.059, 
    353.9068, 353.1668, 353.0458, 352.5217, 352.3766, 351.9774, 351.6346, 
    351.9486, 352.2658, 353.1674, 353.9791, 354.8638, 355.0805, 356.1119, 
    355.2715, 356.6572, 355.4779, 357.5194, 353.8513, 355.4444, 352.5581, 
    352.8694, 353.4318, 354.7221, 354.0263, 354.8403, 353.0411, 352.1061, 
    351.8531, 351.4018, 351.8634, 351.8259, 352.2794, 352.1375, 353.1973, 
    352.6281, 354.2447, 354.834, 356.498, 357.5168, 358.5541, 359.0115, 
    359.1507, 359.2089 ;

 FSH_G =
  354.6916, 355.6444, 355.4608, 356.2226, 355.8003, 356.2989, 354.8835, 
    355.6817, 355.1696, 354.7771, 357.6992, 356.2567, 359.211, 358.2796, 
    360.6015, 359.0676, 360.9107, 360.5579, 361.6212, 361.3167, 362.6746, 
    361.7617, 363.379, 362.457, 362.601, 361.7315, 356.5477, 357.5195, 
    356.4899, 356.6286, 356.5665, 355.8088, 355.4265, 354.6198, 354.765, 
    355.3597, 356.6909, 356.2396, 357.3781, 357.3524, 358.6188, 358.0479, 
    360.1874, 359.5831, 361.3294, 360.8903, 361.3087, 361.1819, 361.3103, 
    360.6663, 360.9422, 360.3756, 358.1547, 358.8158, 356.8665, 355.6996, 
    354.9181, 354.3683, 354.446, 354.5941, 355.3632, 356.0793, 356.6248, 
    356.9894, 357.3488, 358.4343, 359.0219, 360.3093, 360.0776, 360.4706, 
    360.8466, 361.4771, 361.3735, 361.6511, 360.4606, 361.2517, 359.9454, 
    360.3027, 357.4443, 356.3615, 355.8992, 355.4961, 354.5057, 355.1843, 
    354.9167, 355.5612, 355.9655, 355.7656, 356.9994, 356.5197, 359.056, 
    357.9572, 360.8028, 360.1252, 360.9652, 360.5367, 361.2707, 360.6102, 
    361.7545, 362.0034, 361.8333, 362.4873, 360.5735, 361.3085, 355.7599, 
    355.7925, 355.9445, 355.2762, 355.2277, 354.6157, 355.1605, 355.3999, 
    355.9891, 356.3371, 356.668, 357.3953, 358.2069, 359.3537, 360.1691, 
    360.7153, 360.3805, 360.6761, 360.3456, 360.1908, 361.91, 360.9447, 
    362.3932, 362.3132, 361.6576, 362.3222, 355.8154, 355.6279, 354.9682, 
    355.4861, 354.549, 355.0691, 355.3755, 356.5293, 356.7832, 357.018, 
    357.482, 358.0771, 359.1323, 360.0401, 360.8686, 360.808, 360.8293, 
    361.0141, 360.556, 361.0893, 361.1786, 360.9448, 362.3025, 361.9147, 
    362.3115, 362.0591, 355.6889, 356.0045, 355.834, 356.1546, 355.9286, 
    356.933, 357.2341, 358.6427, 358.0653, 358.9966, 358.1589, 358.3051, 
    359.0258, 358.2037, 359.9896, 358.7862, 361.0213, 359.8194, 361.0965, 
    360.865, 361.2485, 361.5917, 362.0237, 362.8199, 362.6356, 363.3015, 
    356.4753, 356.8843, 356.8487, 357.277, 357.5936, 358.2801, 359.392, 
    358.9785, 359.738, 359.8903, 358.7366, 359.4447, 357.1584, 357.5256, 
    357.3073, 356.5073, 359.0732, 357.7509, 360.1825, 359.4731, 361.5427, 
    360.5134, 362.5341, 363.3961, 364.2088, 365.1558, 357.108, 356.83, 
    357.328, 358.0161, 358.6672, 359.5163, 359.6034, 359.7622, 360.1742, 
    360.5204, 359.8121, 360.6071, 357.61, 359.1871, 356.7245, 357.4623, 
    357.9757, 357.7509, 358.9313, 359.2065, 360.3242, 359.7468, 363.183, 
    361.6636, 365.8778, 364.701, 356.7328, 357.1072, 358.4091, 357.7898, 
    359.5732, 360.0088, 360.3632, 360.8155, 360.8646, 361.1325, 360.6934, 
    361.1153, 359.5181, 360.2321, 358.2608, 358.7495, 358.5184, 358.2776, 
    359.0325, 359.8232, 359.8407, 360.094, 360.8065, 359.5804, 363.3778, 
    361.0326, 357.5154, 358.2353, 358.3388, 358.0599, 359.9651, 359.2792, 
    361.1261, 360.6273, 361.4447, 361.0385, 360.9787, 360.457, 360.1319, 
    359.3105, 358.6303, 358.1004, 358.2237, 358.8175, 359.8716, 360.8687, 
    360.6503, 361.3826, 359.4447, 360.2573, 359.9431, 360.7623, 358.9674, 
    360.494, 358.5649, 358.745, 359.2656, 360.3119, 360.5443, 360.7912, 
    360.6389, 359.8985, 359.7775, 359.2531, 359.1079, 358.7084, 358.3655, 
    358.6797, 358.997, 359.8991, 360.7112, 361.5965, 361.8133, 362.8452, 
    362.0043, 363.3908, 362.2108, 364.2535, 360.5834, 362.1774, 359.2895, 
    359.601, 360.1636, 361.4547, 360.7585, 361.5729, 359.7728, 358.8372, 
    358.5841, 358.1325, 358.5945, 358.5569, 359.0107, 358.8687, 359.929, 
    359.3596, 360.977, 361.5667, 363.2316, 364.2509, 365.2888, 365.7464, 
    365.8857, 365.9439 ;

 FSH_NODYNLNDUSE =
  347.9627, 348.915, 348.7315, 349.4929, 349.0708, 349.5691, 348.1545, 
    348.9522, 348.4404, 348.0481, 350.9688, 349.5269, 352.4797, 351.5487, 
    353.8694, 352.3363, 354.1785, 353.8258, 354.8885, 354.5842, 355.9413, 
    355.029, 356.6454, 355.7238, 355.8678, 354.9987, 349.8177, 350.7891, 
    349.76, 349.8986, 349.8366, 349.0793, 348.6972, 347.8909, 348.036, 
    348.6305, 349.961, 349.5098, 350.6478, 350.6221, 351.8878, 351.3172, 
    353.4556, 352.8515, 354.5969, 354.1581, 354.5762, 354.4495, 354.5778, 
    353.9342, 354.21, 353.6437, 351.424, 352.0847, 350.1364, 348.9702, 
    348.1891, 347.6396, 347.7173, 347.8652, 348.6339, 349.3497, 349.8948, 
    350.2593, 350.6184, 351.7034, 352.2906, 353.5774, 353.3458, 353.7385, 
    354.1144, 354.7446, 354.641, 354.9184, 353.7285, 354.5192, 353.2137, 
    353.5708, 350.714, 349.6317, 349.1696, 348.7667, 347.7769, 348.4551, 
    348.1878, 348.8318, 349.2359, 349.0362, 350.2693, 349.7899, 352.3247, 
    351.2266, 354.0706, 353.3933, 354.2329, 353.8047, 354.5382, 353.8781, 
    355.0218, 355.2705, 355.1005, 355.7542, 353.8414, 354.576, 349.0305, 
    349.063, 349.215, 348.5469, 348.4986, 347.8868, 348.4313, 348.6707, 
    349.2595, 349.6073, 349.938, 350.6649, 351.4761, 352.6223, 353.4372, 
    353.9831, 353.6486, 353.9439, 353.6136, 353.4589, 355.1772, 354.2124, 
    355.6602, 355.5802, 354.9249, 355.5892, 349.0859, 348.8985, 348.2392, 
    348.7568, 347.8202, 348.34, 348.6463, 349.7994, 350.0532, 350.2878, 
    350.7516, 351.3464, 352.401, 353.3083, 354.1364, 354.0757, 354.097, 
    354.2818, 353.8239, 354.357, 354.4462, 354.2125, 355.5694, 355.1819, 
    355.5785, 355.3262, 348.9595, 349.275, 349.1045, 349.425, 349.199, 
    350.2029, 350.5038, 351.9117, 351.3346, 352.2654, 351.4281, 351.5743, 
    352.2945, 351.4729, 353.2579, 352.0551, 354.2889, 353.0877, 354.3642, 
    354.1328, 354.5161, 354.859, 355.2908, 356.0865, 355.9024, 356.568, 
    349.7454, 350.1542, 350.1187, 350.5467, 350.8631, 351.5492, 352.6606, 
    352.2473, 353.0063, 353.1586, 352.0056, 352.7132, 350.4281, 350.7952, 
    350.5769, 349.7774, 352.342, 351.0203, 353.4506, 352.7416, 354.8101, 
    353.7813, 355.8009, 356.6625, 357.4747, 358.4212, 350.3778, 350.1, 
    350.5977, 351.2854, 351.9362, 352.7848, 352.8718, 353.0306, 353.4424, 
    353.7883, 353.0804, 353.875, 350.8795, 352.4558, 349.9946, 350.732, 
    351.2451, 351.0204, 352.2001, 352.4752, 353.5923, 353.0151, 356.4496, 
    354.9309, 359.1428, 357.9667, 350.0028, 350.377, 351.6782, 351.0593, 
    352.8416, 353.277, 353.6312, 354.0833, 354.1323, 354.4001, 353.9612, 
    354.3829, 352.7866, 353.5002, 351.53, 352.0184, 351.7875, 351.5468, 
    352.3012, 353.0915, 353.109, 353.3622, 354.0744, 352.8488, 356.6443, 
    354.3003, 350.7849, 351.5045, 351.608, 351.3292, 353.2333, 352.5478, 
    354.3937, 353.8951, 354.7121, 354.3062, 354.2464, 353.7249, 353.4001, 
    352.5791, 351.8992, 351.3697, 351.4929, 352.0864, 353.14, 354.1365, 
    353.9182, 354.65, 352.7133, 353.5253, 353.2113, 354.0301, 352.2362, 
    353.762, 351.8339, 352.0139, 352.5342, 353.58, 353.8122, 354.059, 
    353.9068, 353.1668, 353.0458, 352.5217, 352.3766, 351.9774, 351.6346, 
    351.9486, 352.2658, 353.1674, 353.9791, 354.8638, 355.0805, 356.1119, 
    355.2715, 356.6572, 355.4779, 357.5194, 353.8513, 355.4444, 352.5581, 
    352.8694, 353.4318, 354.7221, 354.0263, 354.8403, 353.0411, 352.1061, 
    351.8531, 351.4018, 351.8634, 351.8259, 352.2794, 352.1375, 353.1973, 
    352.6281, 354.2447, 354.834, 356.498, 357.5168, 358.5541, 359.0115, 
    359.1507, 359.2089 ;

 FSH_R =
  347.9627, 348.915, 348.7315, 349.4929, 349.0708, 349.5691, 348.1545, 
    348.9522, 348.4404, 348.0481, 350.9688, 349.5269, 352.4797, 351.5487, 
    353.8694, 352.3363, 354.1785, 353.8258, 354.8885, 354.5842, 355.9413, 
    355.029, 356.6454, 355.7238, 355.8678, 354.9987, 349.8177, 350.7891, 
    349.76, 349.8986, 349.8366, 349.0793, 348.6972, 347.8909, 348.036, 
    348.6305, 349.961, 349.5098, 350.6478, 350.6221, 351.8878, 351.3172, 
    353.4556, 352.8515, 354.5969, 354.1581, 354.5762, 354.4495, 354.5778, 
    353.9342, 354.21, 353.6437, 351.424, 352.0847, 350.1364, 348.9702, 
    348.1891, 347.6396, 347.7173, 347.8652, 348.6339, 349.3497, 349.8948, 
    350.2593, 350.6184, 351.7034, 352.2906, 353.5774, 353.3458, 353.7385, 
    354.1144, 354.7446, 354.641, 354.9184, 353.7285, 354.5192, 353.2137, 
    353.5708, 350.714, 349.6317, 349.1696, 348.7667, 347.7769, 348.4551, 
    348.1878, 348.8318, 349.2359, 349.0362, 350.2693, 349.7899, 352.3247, 
    351.2266, 354.0706, 353.3933, 354.2329, 353.8047, 354.5382, 353.8781, 
    355.0218, 355.2705, 355.1005, 355.7542, 353.8414, 354.576, 349.0305, 
    349.063, 349.215, 348.5469, 348.4986, 347.8868, 348.4313, 348.6707, 
    349.2595, 349.6073, 349.938, 350.6649, 351.4761, 352.6223, 353.4372, 
    353.9831, 353.6486, 353.9439, 353.6136, 353.4589, 355.1772, 354.2124, 
    355.6602, 355.5802, 354.9249, 355.5892, 349.0859, 348.8985, 348.2392, 
    348.7568, 347.8202, 348.34, 348.6463, 349.7994, 350.0532, 350.2878, 
    350.7516, 351.3464, 352.401, 353.3083, 354.1364, 354.0757, 354.097, 
    354.2818, 353.8239, 354.357, 354.4462, 354.2125, 355.5694, 355.1819, 
    355.5785, 355.3262, 348.9595, 349.275, 349.1045, 349.425, 349.199, 
    350.2029, 350.5038, 351.9117, 351.3346, 352.2654, 351.4281, 351.5743, 
    352.2945, 351.4729, 353.2579, 352.0551, 354.2889, 353.0877, 354.3642, 
    354.1328, 354.5161, 354.859, 355.2908, 356.0865, 355.9024, 356.568, 
    349.7454, 350.1542, 350.1187, 350.5467, 350.8631, 351.5492, 352.6606, 
    352.2473, 353.0063, 353.1586, 352.0056, 352.7132, 350.4281, 350.7952, 
    350.5769, 349.7774, 352.342, 351.0203, 353.4506, 352.7416, 354.8101, 
    353.7813, 355.8009, 356.6625, 357.4747, 358.4212, 350.3778, 350.1, 
    350.5977, 351.2854, 351.9362, 352.7848, 352.8718, 353.0306, 353.4424, 
    353.7883, 353.0804, 353.875, 350.8795, 352.4558, 349.9946, 350.732, 
    351.2451, 351.0204, 352.2001, 352.4752, 353.5923, 353.0151, 356.4496, 
    354.9309, 359.1428, 357.9667, 350.0028, 350.377, 351.6782, 351.0593, 
    352.8416, 353.277, 353.6312, 354.0833, 354.1323, 354.4001, 353.9612, 
    354.3829, 352.7866, 353.5002, 351.53, 352.0184, 351.7875, 351.5468, 
    352.3012, 353.0915, 353.109, 353.3622, 354.0744, 352.8488, 356.6443, 
    354.3003, 350.7849, 351.5045, 351.608, 351.3292, 353.2333, 352.5478, 
    354.3937, 353.8951, 354.7121, 354.3062, 354.2464, 353.7249, 353.4001, 
    352.5791, 351.8992, 351.3697, 351.4929, 352.0864, 353.14, 354.1365, 
    353.9182, 354.65, 352.7133, 353.5253, 353.2113, 354.0301, 352.2362, 
    353.762, 351.8339, 352.0139, 352.5342, 353.58, 353.8122, 354.059, 
    353.9068, 353.1668, 353.0458, 352.5217, 352.3766, 351.9774, 351.6346, 
    351.9486, 352.2658, 353.1674, 353.9791, 354.8638, 355.0805, 356.1119, 
    355.2715, 356.6572, 355.4779, 357.5194, 353.8513, 355.4444, 352.5581, 
    352.8694, 353.4318, 354.7221, 354.0263, 354.8403, 353.0411, 352.1061, 
    351.8531, 351.4018, 351.8634, 351.8259, 352.2794, 352.1375, 353.1973, 
    352.6281, 354.2447, 354.834, 356.498, 357.5168, 358.5541, 359.0115, 
    359.1507, 359.2089 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.728875, -6.729403, -6.729306, -6.729714, -6.729492, -6.729756, 
    -6.728984, -6.729419, -6.729139, -6.728928, -6.730493, -6.729734, 
    -6.731331, -6.730838, -6.732092, -6.731248, -6.732265, -6.73208, 
    -6.732666, -6.732499, -6.733226, -6.732744, -6.733623, -6.733117, 
    -6.733192, -6.732726, -6.729897, -6.730395, -6.729865, -6.729937, 
    -6.729907, -6.729493, -6.729277, -6.728844, -6.728922, -6.729248, 
    -6.72997, -6.729732, -6.730353, -6.730339, -6.731024, -6.730715, 
    -6.731876, -6.731549, -6.732506, -6.732263, -6.732492, -6.732425, 
    -6.732493, -6.732138, -6.73229, -6.731981, -6.730771, -6.731122, 
    -6.730068, -6.729419, -6.729001, -6.728706, -6.728748, -6.728825, 
    -6.729249, -6.729644, -6.729942, -6.73014, -6.730337, -6.730903, 
    -6.731228, -6.731937, -6.731819, -6.732027, -6.73224, -6.732584, 
    -6.732529, -6.732678, -6.732028, -6.732457, -6.731749, -6.731941, 
    -6.730352, -6.729797, -6.729529, -6.729323, -6.728779, -6.729143, 
    -6.728998, -6.729364, -6.729582, -6.729476, -6.730146, -6.729884, 
    -6.731247, -6.730659, -6.732215, -6.731844, -6.732305, -6.732071, 
    -6.732469, -6.732111, -6.732737, -6.732869, -6.732778, -6.733141, 
    -6.73209, -6.732489, -6.729471, -6.729488, -6.729572, -6.729202, 
    -6.729167, -6.72884, -6.729135, -6.729272, -6.729598, -6.729784, 
    -6.729963, -6.730358, -6.730794, -6.731415, -6.731867, -6.732169, 
    -6.731987, -6.732148, -6.731966, -6.731883, -6.732817, -6.732289, 
    -6.733088, -6.733046, -6.73268, -6.73305, -6.729501, -6.729402, 
    -6.729029, -6.729324, -6.728805, -6.729082, -6.729254, -6.729881, 
    -6.730028, -6.730153, -6.730408, -6.73073, -6.731296, -6.731793, 
    -6.732254, -6.732221, -6.732232, -6.732331, -6.73208, -6.732372, 
    -6.732418, -6.732294, -6.733039, -6.732827, -6.733045, -6.732907, 
    -6.729435, -6.729604, -6.729512, -6.729683, -6.729559, -6.730098, 
    -6.73026, -6.731028, -6.730722, -6.73122, -6.730775, -6.730852, -6.73122, 
    -6.730802, -6.731758, -6.731096, -6.732335, -6.731657, -6.732377, 
    -6.732252, -6.732462, -6.732646, -6.732886, -6.733317, -6.733219, 
    -6.733586, -6.72986, -6.730076, -6.730064, -6.730296, -6.730465, 
    -6.730843, -6.731441, -6.731218, -6.731634, -6.731715, -6.731087, 
    -6.731466, -6.730227, -6.730419, -6.73031, -6.729873, -6.731259, 
    -6.730543, -6.731874, -6.731486, -6.732619, -6.732048, -6.733163, 
    -6.733622, -6.734088, -6.734595, -6.730202, -6.730054, -6.730326, 
    -6.730688, -6.731045, -6.731509, -6.73156, -6.731645, -6.731874, 
    -6.732062, -6.731665, -6.73211, -6.730449, -6.731325, -6.729992, 
    -6.730383, -6.730669, -6.730551, -6.731194, -6.731344, -6.731947, 
    -6.731639, -6.733502, -6.732676, -6.735005, -6.734348, -6.730001, 
    -6.730205, -6.730906, -6.730573, -6.731544, -6.731779, -6.731977, 
    -6.732219, -6.73225, -6.732394, -6.732157, -6.732388, -6.73151, 
    -6.731903, -6.730834, -6.73109, -6.730975, -6.730843, -6.731249, 
    -6.731669, -6.731689, -6.731822, -6.732177, -6.731548, -6.733588, 
    -6.732306, -6.730427, -6.730805, -6.730873, -6.730724, -6.731755, 
    -6.73138, -6.732392, -6.732121, -6.732569, -6.732345, -6.732312, 
    -6.732028, -6.731847, -6.731395, -6.73103, -6.730747, -6.730814, 
    -6.731125, -6.731698, -6.732248, -6.732126, -6.732535, -6.731472, 
    -6.731912, -6.731738, -6.732193, -6.73121, -6.732012, -6.731, -6.731091, 
    -6.731373, -6.731934, -6.732075, -6.732205, -6.732127, -6.731714, 
    -6.731652, -6.731369, -6.731285, -6.731073, -6.730891, -6.731054, 
    -6.731223, -6.731719, -6.732161, -6.732647, -6.732771, -6.733312, 
    -6.732856, -6.733593, -6.732942, -6.734081, -6.732075, -6.732946, 
    -6.73139, -6.731559, -6.731855, -6.732559, -6.732191, -6.732627, 
    -6.73165, -6.73113, -6.731009, -6.730762, -6.731015, -6.730995, 
    -6.731237, -6.731161, -6.731736, -6.731427, -6.732308, -6.732626, 
    -6.733543, -6.734099, -6.734684, -6.734937, -6.735015, -6.735047 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  2.413656e-36, 2.065401e-35, 1.367197e-35, 7.458777e-35, 2.924233e-35, 
    8.819833e-35, 3.748208e-36, 2.246482e-35, 7.197595e-36, 2.935293e-36, 
    1.796957e-33, 8.037766e-35, 3.922441e-32, 6.007093e-33, 6.052333e-31, 
    2.939911e-32, 1.094422e-30, 5.556852e-31, 4.175555e-30, 2.359349e-30, 
    2.893847e-29, 5.424175e-30, 1.017046e-28, 1.948533e-29, 2.531664e-29, 
    5.128552e-30, 1.5186e-34, 1.229759e-33, 1.339012e-34, 1.812237e-34, 
    1.582295e-34, 2.981927e-35, 1.267358e-35, 2.04289e-36, 2.854736e-36, 
    1.088977e-35, 2.075535e-34, 7.733206e-35, 9.06774e-34, 8.585492e-34, 
    1.206895e-32, 3.712564e-33, 2.708682e-31, 8.236855e-32, 2.416494e-30, 
    1.051322e-30, 2.324528e-30, 1.82943e-30, 2.331775e-30, 6.847458e-31, 
    1.161084e-30, 3.905416e-31, 4.637344e-33, 1.761981e-32, 3.033677e-34, 
    2.342121e-35, 4.05827e-36, 1.140883e-36, 1.366814e-36, 1.926661e-36, 
    1.097471e-35, 5.431533e-35, 1.795261e-34, 3.950291e-34, 8.518304e-34, 
    8.288211e-33, 2.678748e-32, 3.436761e-31, 2.184636e-31, 4.697071e-31, 
    9.671604e-31, 3.190841e-30, 2.625917e-30, 4.41738e-30, 4.603185e-31, 
    2.088884e-30, 1.685259e-31, 3.389846e-31, 1.048926e-33, 1.010662e-34, 
    3.652738e-35, 1.480341e-35, 1.570089e-36, 7.446789e-36, 4.047018e-36, 
    1.712407e-35, 4.221452e-35, 2.705511e-35, 4.035902e-34, 1.42863e-34, 
    2.869719e-32, 3.075397e-33, 8.894096e-31, 2.398156e-31, 1.212633e-30, 
    5.331979e-31, 2.164703e-30, 6.143018e-31, 5.354316e-30, 8.491746e-30, 
    6.198718e-30, 2.057202e-29, 5.724397e-31, 2.324658e-30, 2.671984e-35, 
    2.873639e-35, 4.028986e-35, 9.014748e-36, 8.217192e-36, 2.024267e-36, 
    7.050135e-36, 1.192036e-35, 4.446345e-35, 9.581258e-35, 1.972759e-34, 
    9.40965e-34, 5.171452e-33, 5.218879e-32, 2.613056e-31, 7.518973e-31, 
    3.941118e-31, 6.973537e-31, 3.683514e-31, 2.724792e-31, 7.147453e-30, 
    1.166841e-30, 1.73386e-29, 1.498157e-29, 4.472238e-30, 1.523048e-29, 
    3.024102e-35, 1.988205e-35, 4.550449e-36, 1.44646e-35, 1.73507e-36, 
    5.729078e-36, 1.12904e-35, 1.460426e-34, 2.53197e-34, 4.202358e-34, 
    1.130701e-33, 3.94548e-33, 3.344858e-32, 2.031258e-31, 1.00837e-30, 
    8.979328e-31, 9.353917e-31, 1.33104e-30, 5.534872e-31, 1.535411e-30, 
    1.819247e-30, 1.166494e-30, 1.469084e-29, 7.203947e-30, 1.493503e-29, 
    9.401376e-30, 2.279148e-35, 4.603192e-35, 3.151121e-35, 6.416304e-35, 
    3.891003e-35, 3.504587e-34, 6.685744e-34, 1.269163e-32, 3.850616e-33, 
    2.54377e-32, 4.67595e-33, 6.33306e-33, 2.703684e-32, 5.129652e-33, 
    1.84164e-31, 1.661233e-32, 1.349351e-30, 1.31887e-31, 1.556519e-30, 
    1.001499e-30, 2.074591e-30, 3.953509e-30, 8.809192e-30, 3.754736e-29, 
    2.692728e-29, 8.862534e-29, 1.296324e-34, 3.153121e-34, 2.916695e-34, 
    7.313115e-34, 1.432144e-33, 6.009421e-33, 5.630612e-32, 2.449265e-32, 
    1.119704e-31, 1.512694e-31, 1.497909e-32, 6.257924e-32, 5.680003e-34, 
    1.242106e-33, 7.802933e-34, 1.391165e-34, 2.970523e-32, 1.996976e-33, 
    2.682689e-31, 6.618635e-32, 3.607827e-30, 5.103762e-31, 2.240553e-29, 
    1.049413e-28, 4.315611e-28, 2.151595e-27, 5.097033e-34, 2.801228e-34, 
    8.151042e-34, 3.479038e-33, 1.300711e-32, 7.215027e-32, 8.574919e-32, 
    1.175121e-31, 2.638394e-31, 5.166526e-31, 1.297972e-31, 6.107406e-31, 
    1.487772e-33, 3.735418e-32, 2.231189e-34, 1.086605e-33, 3.196354e-33, 
    1.995071e-33, 2.225378e-32, 3.879716e-32, 3.537037e-31, 1.139286e-31, 
    7.1979e-29, 4.527107e-30, 7.072285e-27, 1.001204e-27, 2.26989e-34, 
    5.086269e-34, 7.850772e-33, 2.164587e-33, 8.075713e-32, 1.909646e-31, 
    3.810726e-31, 9.116114e-31, 1.000794e-30, 1.666826e-30, 7.208881e-31, 
    1.612822e-30, 7.241077e-32, 2.954449e-31, 5.773067e-33, 1.538488e-32, 
    9.818068e-33, 5.978102e-33, 2.731482e-32, 1.326861e-31, 1.371577e-31, 
    2.257592e-31, 9.004322e-31, 8.191729e-32, 1.019036e-28, 1.384652e-30, 
    1.213156e-33, 5.487309e-33, 6.787049e-33, 3.804815e-33, 1.752723e-31, 
    4.491113e-32, 1.646268e-30, 6.348694e-31, 3.001185e-30, 1.393988e-30, 
    1.244232e-30, 4.570806e-31, 2.430007e-31, 4.783712e-32, 1.235653e-32, 
    4.139165e-33, 5.346258e-33, 1.767639e-32, 1.459641e-31, 1.009369e-30, 
    6.642821e-31, 2.670752e-30, 6.253374e-32, 3.104628e-31, 1.679492e-31, 
    8.230366e-31, 2.39545e-32, 4.932957e-31, 1.079973e-32, 1.5238e-32, 
    4.370052e-32, 3.45641e-31, 5.410543e-31, 8.702187e-31, 6.493018e-31, 
    1.538556e-31, 1.211231e-31, 4.260206e-32, 3.183188e-32, 1.413956e-32, 
    7.167403e-33, 1.333833e-32, 2.544929e-32, 1.539362e-31, 7.466343e-31, 
    3.989861e-30, 5.969769e-30, 3.938643e-29, 8.521178e-30, 1.042838e-28, 
    1.24947e-29, 4.677264e-28, 5.850539e-31, 1.171975e-29, 4.582477e-32, 
    8.533778e-32, 2.588349e-31, 3.063866e-30, 8.169875e-31, 3.821891e-30, 
    1.199891e-31, 1.841584e-32, 1.123526e-32, 4.426199e-33, 1.147535e-32, 
    1.062511e-32, 2.613189e-32, 1.959549e-32, 1.632738e-31, 5.273784e-32, 
    1.240751e-30, 3.776026e-30, 7.832231e-29, 4.6458e-28, 2.680098e-27, 
    5.702732e-27, 7.160027e-27, 7.872312e-27 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1.95279e-35, 1.671031e-34, 1.106143e-34, 6.034591e-34, 2.365878e-34, 
    7.135766e-34, 3.032522e-35, 1.817537e-34, 5.823279e-35, 2.374826e-35, 
    1.453844e-32, 6.503028e-34, 3.173486e-31, 4.860093e-32, 4.896695e-30, 
    2.378562e-31, 8.854517e-30, 4.495822e-30, 3.378271e-29, 1.908853e-29, 
    2.341293e-28, 4.388478e-29, 8.228507e-28, 1.576479e-28, 2.048266e-28, 
    4.149302e-29, 1.228637e-33, 9.949474e-33, 1.08334e-33, 1.466207e-33, 
    1.28017e-33, 2.412555e-34, 1.025367e-34, 1.652819e-35, 2.30965e-35, 
    8.810464e-35, 1.679231e-33, 6.256621e-34, 7.336337e-33, 6.94617e-33, 
    9.76449e-32, 3.003683e-32, 2.191484e-30, 6.664103e-31, 1.955087e-29, 
    8.505818e-30, 1.880681e-29, 1.480117e-29, 1.886544e-29, 5.539998e-30, 
    9.393852e-30, 3.159713e-30, 3.751885e-32, 1.425547e-31, 2.454424e-33, 
    1.894914e-34, 3.283381e-35, 9.230414e-36, 1.105833e-35, 1.558783e-35, 
    8.879191e-35, 4.394431e-34, 1.452472e-33, 3.196019e-33, 6.891812e-33, 
    6.705652e-32, 2.167266e-31, 2.780543e-30, 1.767499e-30, 3.800208e-30, 
    7.824898e-30, 2.581579e-29, 2.124522e-29, 3.573922e-29, 3.724249e-30, 
    1.690031e-29, 1.363474e-30, 2.742586e-30, 8.486433e-33, 8.176849e-34, 
    2.955281e-34, 1.197683e-34, 1.270295e-35, 6.024892e-35, 3.274277e-35, 
    1.385438e-34, 3.415405e-34, 2.188918e-34, 3.265283e-33, 1.155846e-33, 
    2.321772e-31, 2.488178e-32, 7.195849e-30, 1.94025e-30, 9.810919e-30, 
    4.313886e-30, 1.751373e-29, 4.970064e-30, 4.331958e-29, 6.870325e-29, 
    5.01513e-29, 1.664398e-28, 4.631375e-30, 1.880786e-29, 2.161793e-34, 
    2.324944e-34, 3.259688e-34, 7.293464e-35, 6.648194e-35, 1.637752e-35, 
    5.703976e-35, 9.644278e-35, 3.597356e-34, 7.751804e-34, 1.596078e-33, 
    7.612963e-33, 4.184011e-32, 4.222381e-31, 2.114117e-30, 6.083293e-30, 
    3.188597e-30, 5.642004e-30, 2.98018e-30, 2.204518e-30, 5.782712e-29, 
    9.440435e-30, 1.402795e-28, 1.212097e-28, 3.618305e-29, 1.232236e-28, 
    2.446677e-34, 1.608575e-34, 3.681582e-35, 1.170272e-34, 1.403774e-35, 
    4.635162e-35, 9.134602e-35, 1.181571e-33, 2.048513e-33, 3.399956e-33, 
    9.148041e-33, 3.192127e-32, 2.706188e-31, 1.643407e-30, 8.158312e-30, 
    7.264806e-30, 7.567872e-30, 1.07689e-29, 4.478038e-30, 1.242238e-29, 
    1.471879e-29, 9.437629e-30, 1.188575e-28, 5.828419e-29, 1.208332e-28, 
    7.606269e-29, 1.843965e-34, 3.724254e-34, 2.549443e-34, 5.191169e-34, 
    3.148051e-34, 2.835418e-33, 5.409163e-33, 1.026828e-31, 3.115376e-32, 
    2.058061e-31, 3.78312e-32, 5.123819e-32, 2.18744e-31, 4.150192e-32, 
    1.489996e-30, 1.344036e-31, 1.091705e-29, 1.067044e-30, 1.259316e-29, 
    8.102715e-30, 1.678467e-29, 3.198622e-29, 7.127157e-29, 3.037804e-28, 
    2.178576e-28, 7.170314e-28, 1.048803e-33, 2.551061e-33, 2.359779e-33, 
    5.916742e-33, 1.158689e-32, 4.861977e-32, 4.555498e-31, 1.9816e-31, 
    9.059063e-31, 1.223859e-30, 1.211897e-31, 5.06303e-31, 4.595458e-33, 
    1.004937e-32, 6.313034e-33, 1.125535e-33, 2.403329e-31, 1.615672e-32, 
    2.170454e-30, 5.354867e-31, 2.918945e-29, 4.129245e-30, 1.812739e-28, 
    8.490375e-28, 3.491585e-27, 1.740767e-26, 4.123801e-33, 2.266359e-33, 
    6.594675e-33, 2.814747e-32, 1.052352e-31, 5.837384e-31, 6.937616e-31, 
    9.50742e-31, 2.134617e-30, 4.180025e-30, 1.050136e-30, 4.941253e-30, 
    1.203695e-32, 3.022174e-31, 1.805164e-33, 8.791276e-33, 2.586039e-32, 
    1.614131e-32, 1.800462e-31, 3.138919e-31, 2.861672e-30, 9.217499e-31, 
    5.823526e-28, 3.662697e-29, 5.721897e-26, 8.100334e-27, 1.836475e-33, 
    4.115093e-33, 6.351738e-32, 1.751279e-32, 6.533729e-31, 1.545017e-30, 
    3.083102e-30, 7.375475e-30, 8.097016e-30, 1.348561e-29, 5.832411e-30, 
    1.304868e-29, 5.858459e-31, 2.390324e-30, 4.670752e-32, 1.244728e-31, 
    7.943397e-32, 4.836638e-32, 2.20993e-31, 1.073509e-30, 1.109687e-30, 
    1.826525e-30, 7.285029e-30, 6.627593e-31, 8.244606e-28, 1.120265e-29, 
    9.815149e-33, 4.439557e-32, 5.491123e-32, 3.078321e-32, 1.418056e-30, 
    3.633576e-31, 1.331928e-29, 5.136468e-30, 2.428136e-29, 1.127819e-29, 
    1.006657e-29, 3.698052e-30, 1.966019e-30, 3.870306e-31, 9.997165e-32, 
    3.348829e-32, 4.325439e-32, 1.430124e-31, 1.180936e-30, 8.166389e-30, 
    5.374434e-30, 2.160796e-29, 5.059349e-31, 2.511828e-30, 1.358808e-30, 
    6.658852e-30, 1.938061e-31, 3.991053e-30, 8.737623e-32, 1.232844e-31, 
    3.535631e-31, 2.79644e-30, 4.377449e-30, 7.040583e-30, 5.253235e-30, 
    1.244783e-30, 9.799575e-31, 3.446758e-31, 2.575388e-31, 1.143974e-31, 
    5.798853e-32, 1.07915e-31, 2.058998e-31, 1.245435e-30, 6.040713e-30, 
    3.228034e-29, 4.829896e-29, 3.186595e-28, 6.894137e-29, 8.437176e-28, 
    1.010895e-28, 3.784183e-27, 4.733432e-30, 9.481973e-29, 3.707495e-31, 
    6.904331e-31, 2.094127e-30, 2.478849e-29, 6.609912e-30, 3.092136e-29, 
    9.707829e-31, 1.489951e-31, 9.08999e-32, 3.581057e-32, 9.284234e-32, 
    8.596343e-32, 2.114224e-31, 1.585391e-31, 1.320982e-30, 4.266803e-31, 
    1.003841e-29, 3.055028e-29, 6.336738e-28, 3.758727e-27, 2.168357e-26, 
    4.613847e-26, 5.792885e-26, 6.369166e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  5.215076e-38, 4.462618e-37, 2.954041e-37, 1.611585e-36, 6.318259e-37, 
    1.905662e-36, 8.098581e-38, 4.853872e-37, 1.555152e-37, 6.342154e-38, 
    3.882606e-35, 1.736684e-36, 8.475047e-34, 1.297926e-34, 1.307701e-32, 
    6.352137e-34, 2.364669e-32, 1.200645e-32, 9.02194e-32, 5.097743e-32, 
    6.252607e-31, 1.171978e-31, 2.197487e-30, 4.21011e-31, 5.470054e-31, 
    1.108104e-31, 3.281171e-36, 2.657085e-35, 2.893143e-36, 3.915621e-36, 
    3.418794e-36, 6.442916e-37, 2.738322e-37, 4.413979e-38, 6.168097e-38, 
    2.352902e-37, 4.484517e-36, 1.670879e-36, 1.959227e-35, 1.855029e-35, 
    2.607684e-34, 8.021573e-35, 5.852531e-33, 1.779701e-33, 5.221213e-32, 
    2.271546e-32, 5.022506e-32, 3.95277e-32, 5.038164e-32, 1.4795e-32, 
    2.508702e-32, 8.438263e-33, 1.00197e-34, 3.807036e-34, 6.554731e-36, 
    5.060515e-37, 8.768519e-38, 2.465052e-38, 2.953212e-38, 4.162849e-38, 
    2.371256e-37, 1.173567e-36, 3.87894e-36, 8.535219e-36, 1.840512e-35, 
    1.790797e-34, 5.787855e-34, 7.425659e-33, 4.720247e-33, 1.014876e-32, 
    2.089701e-32, 6.894311e-32, 5.673703e-32, 9.544439e-32, 9.945901e-33, 
    4.513361e-32, 3.641265e-33, 7.324293e-33, 2.266369e-35, 2.183691e-36, 
    7.892308e-37, 3.198505e-37, 3.392419e-38, 1.608994e-37, 8.744207e-38, 
    3.69992e-37, 9.121102e-37, 5.845676e-37, 8.720196e-36, 3.086777e-36, 
    6.200476e-34, 6.644875e-35, 1.921708e-32, 5.18159e-33, 2.620083e-32, 
    1.152057e-32, 4.677179e-32, 1.327295e-32, 1.156883e-31, 1.834774e-31, 
    1.33933e-31, 4.444906e-31, 1.236845e-32, 5.022787e-32, 5.773235e-37, 
    6.208942e-37, 8.705248e-37, 1.947776e-37, 1.775451e-37, 4.37374e-38, 
    1.52329e-37, 2.575579e-37, 9.607018e-37, 2.07018e-36, 4.262452e-36, 
    2.033101e-35, 1.117373e-34, 1.12762e-33, 5.645917e-33, 1.624592e-32, 
    8.515401e-33, 1.506742e-32, 7.958807e-33, 5.887339e-33, 1.544319e-31, 
    2.521143e-32, 3.746275e-31, 3.237001e-31, 9.662969e-32, 3.290782e-31, 
    6.534041e-37, 4.295824e-37, 9.831946e-38, 3.125301e-37, 3.748885e-38, 
    1.237856e-37, 2.439466e-37, 3.155478e-36, 5.470714e-36, 9.079849e-36, 
    2.443056e-35, 8.524826e-35, 7.227089e-34, 4.38885e-33, 2.178742e-32, 
    1.940124e-32, 2.02106e-32, 2.87592e-32, 1.195896e-32, 3.317495e-32, 
    3.930768e-32, 2.520394e-32, 3.174184e-31, 1.556525e-31, 3.226945e-31, 
    2.031314e-31, 4.924451e-37, 9.94591e-37, 6.808485e-37, 1.386342e-36, 
    8.407115e-37, 7.572205e-36, 1.444559e-35, 2.742225e-34, 8.319856e-35, 
    5.496213e-34, 1.010312e-34, 1.368356e-34, 5.841733e-34, 1.108341e-34, 
    3.979152e-33, 3.589353e-34, 2.915483e-32, 2.849626e-33, 3.363103e-32, 
    2.163894e-32, 4.482479e-32, 8.542173e-32, 1.903363e-31, 8.112692e-31, 
    5.818058e-31, 1.914888e-30, 2.80091e-36, 6.812808e-36, 6.301973e-36, 
    1.580113e-35, 3.09437e-35, 1.298429e-34, 1.216582e-33, 5.292021e-34, 
    2.419295e-33, 3.268412e-33, 3.236466e-34, 1.352122e-33, 1.227253e-35, 
    2.683763e-35, 1.685945e-35, 3.005829e-36, 6.41828e-34, 4.314779e-35, 
    5.796368e-33, 1.43006e-33, 7.795273e-32, 1.102748e-32, 4.841063e-31, 
    2.26742e-30, 9.324546e-30, 4.648852e-29, 1.101293e-35, 6.052488e-36, 
    1.76116e-35, 7.517005e-35, 2.810389e-34, 1.558919e-33, 1.852745e-33, 
    2.539032e-33, 5.700664e-33, 1.116309e-32, 2.804471e-33, 1.319601e-32, 
    3.214563e-35, 8.070954e-34, 4.820831e-36, 2.347779e-35, 6.906222e-35, 
    4.310663e-35, 4.808277e-34, 8.382732e-34, 7.642322e-33, 2.461606e-33, 
    1.555218e-30, 9.781522e-32, 1.528075e-28, 2.163256e-29, 4.904451e-36, 
    1.098968e-35, 1.696282e-34, 4.676928e-35, 1.744884e-33, 4.126089e-33, 
    8.233669e-33, 1.969679e-32, 2.162372e-32, 3.601439e-32, 1.557591e-32, 
    3.484753e-32, 1.564548e-33, 6.383549e-33, 1.247361e-34, 3.324145e-34, 
    2.121347e-34, 1.291662e-34, 5.901793e-34, 2.86689e-33, 2.963506e-33, 
    4.87788e-33, 1.945524e-32, 1.769951e-33, 2.201786e-30, 2.991757e-32, 
    2.621213e-35, 1.185619e-34, 1.466448e-34, 8.220897e-35, 3.787031e-33, 
    9.703751e-34, 3.55702e-32, 1.371735e-32, 6.484529e-32, 3.01193e-32, 
    2.688357e-32, 9.875941e-33, 5.25041e-33, 1.033596e-33, 2.669822e-34, 
    8.943312e-35, 1.155143e-34, 3.81926e-34, 3.153782e-33, 2.180899e-32, 
    1.435285e-32, 5.770578e-32, 1.351139e-33, 6.708035e-33, 3.628804e-33, 
    1.778299e-32, 5.175745e-34, 1.065842e-32, 2.333451e-34, 3.292408e-34, 
    9.442181e-34, 7.468114e-33, 1.169032e-32, 1.880243e-32, 1.402918e-32, 
    3.324291e-33, 2.617054e-33, 9.204841e-34, 6.877776e-34, 3.055072e-34, 
    1.548629e-34, 2.881955e-34, 5.498716e-34, 3.326032e-33, 1.61322e-32, 
    8.620718e-32, 1.289862e-31, 8.510052e-31, 1.841134e-31, 2.253214e-30, 
    2.699674e-31, 1.010595e-29, 1.2641e-32, 2.532236e-31, 9.901159e-34, 
    1.843856e-33, 5.592533e-33, 6.619962e-32, 1.765229e-32, 8.257793e-32, 
    2.592552e-33, 3.979031e-34, 2.427554e-34, 9.563495e-35, 2.479428e-34, 
    2.295721e-34, 5.646202e-34, 4.233913e-34, 3.527786e-33, 1.139483e-33, 
    2.680836e-32, 8.158694e-32, 1.692275e-30, 1.003797e-29, 5.790762e-29, 
    1.232162e-28, 1.547033e-28, 1.700933e-28 ;

 F_N2O_NIT =
  3.45013e-14, 3.468788e-14, 3.465158e-14, 3.480231e-14, 3.471866e-14, 
    3.481741e-14, 3.453909e-14, 3.469527e-14, 3.459553e-14, 3.451807e-14, 
    3.509563e-14, 3.480903e-14, 3.539461e-14, 3.521096e-14, 3.567316e-14, 
    3.536599e-14, 3.573525e-14, 3.566431e-14, 3.587808e-14, 3.581678e-14, 
    3.609079e-14, 3.590639e-14, 3.623325e-14, 3.604672e-14, 3.607585e-14, 
    3.590029e-14, 3.486666e-14, 3.505991e-14, 3.485522e-14, 3.488274e-14, 
    3.487039e-14, 3.472037e-14, 3.464486e-14, 3.448705e-14, 3.451568e-14, 
    3.46316e-14, 3.48951e-14, 3.480557e-14, 3.503146e-14, 3.502635e-14, 
    3.527859e-14, 3.516476e-14, 3.558998e-14, 3.546888e-14, 3.581933e-14, 
    3.573104e-14, 3.581517e-14, 3.578965e-14, 3.581549e-14, 3.568606e-14, 
    3.574148e-14, 3.562769e-14, 3.518609e-14, 3.531561e-14, 3.492992e-14, 
    3.46989e-14, 3.454591e-14, 3.443752e-14, 3.445283e-14, 3.448203e-14, 
    3.463228e-14, 3.477383e-14, 3.488189e-14, 3.495424e-14, 3.502561e-14, 
    3.524197e-14, 3.53568e-14, 3.561446e-14, 3.556792e-14, 3.56468e-14, 
    3.572226e-14, 3.584908e-14, 3.58282e-14, 3.588412e-14, 3.564472e-14, 
    3.580373e-14, 3.554139e-14, 3.561305e-14, 3.504496e-14, 3.482973e-14, 
    3.473835e-14, 3.465852e-14, 3.44646e-14, 3.459846e-14, 3.454566e-14, 
    3.467134e-14, 3.47513e-14, 3.471174e-14, 3.495622e-14, 3.486107e-14, 
    3.53636e-14, 3.514674e-14, 3.571346e-14, 3.557747e-14, 3.574608e-14, 
    3.566e-14, 3.580754e-14, 3.567474e-14, 3.590494e-14, 3.595515e-14, 
    3.592083e-14, 3.605276e-14, 3.566736e-14, 3.581513e-14, 3.471065e-14, 
    3.47171e-14, 3.474715e-14, 3.461509e-14, 3.460702e-14, 3.448625e-14, 
    3.459371e-14, 3.463951e-14, 3.475594e-14, 3.482487e-14, 3.489046e-14, 
    3.503489e-14, 3.519649e-14, 3.542306e-14, 3.558627e-14, 3.569585e-14, 
    3.562865e-14, 3.568797e-14, 3.562164e-14, 3.559057e-14, 3.593632e-14, 
    3.574198e-14, 3.603376e-14, 3.60176e-14, 3.588542e-14, 3.601941e-14, 
    3.472162e-14, 3.468451e-14, 3.455578e-14, 3.46565e-14, 3.44731e-14, 
    3.457569e-14, 3.463473e-14, 3.486303e-14, 3.491331e-14, 3.495993e-14, 
    3.50521e-14, 3.517055e-14, 3.537879e-14, 3.556043e-14, 3.572664e-14, 
    3.571445e-14, 3.571874e-14, 3.57559e-14, 3.566386e-14, 3.577102e-14, 
    3.578901e-14, 3.574196e-14, 3.601542e-14, 3.59372e-14, 3.601724e-14, 
    3.59663e-14, 3.469657e-14, 3.475903e-14, 3.472526e-14, 3.478875e-14, 
    3.474401e-14, 3.494314e-14, 3.500295e-14, 3.528344e-14, 3.516822e-14, 
    3.535169e-14, 3.518683e-14, 3.521601e-14, 3.535764e-14, 3.519573e-14, 
    3.555038e-14, 3.530973e-14, 3.575734e-14, 3.551635e-14, 3.577246e-14, 
    3.57259e-14, 3.580301e-14, 3.587212e-14, 3.595916e-14, 3.612001e-14, 
    3.608274e-14, 3.621746e-14, 3.485225e-14, 3.493343e-14, 3.49263e-14, 
    3.501135e-14, 3.507431e-14, 3.521098e-14, 3.543067e-14, 3.534799e-14, 
    3.549986e-14, 3.553038e-14, 3.529967e-14, 3.544122e-14, 3.49878e-14, 
    3.506085e-14, 3.501736e-14, 3.48586e-14, 3.536698e-14, 3.510564e-14, 
    3.558893e-14, 3.544684e-14, 3.586225e-14, 3.565536e-14, 3.606222e-14, 
    3.623674e-14, 3.640144e-14, 3.659424e-14, 3.497779e-14, 3.492258e-14, 
    3.502148e-14, 3.515848e-14, 3.528587e-14, 3.545553e-14, 3.547292e-14, 
    3.550474e-14, 3.558726e-14, 3.56567e-14, 3.551478e-14, 3.567411e-14, 
    3.507777e-14, 3.538972e-14, 3.490167e-14, 3.504828e-14, 3.515037e-14, 
    3.510558e-14, 3.533851e-14, 3.53935e-14, 3.561738e-14, 3.550158e-14, 
    3.619361e-14, 3.588668e-14, 3.67414e-14, 3.65016e-14, 3.490329e-14, 
    3.49776e-14, 3.523676e-14, 3.511335e-14, 3.546687e-14, 3.555413e-14, 
    3.562515e-14, 3.571601e-14, 3.572583e-14, 3.577972e-14, 3.569142e-14, 
    3.577623e-14, 3.545586e-14, 3.559886e-14, 3.520708e-14, 3.530225e-14, 
    3.525845e-14, 3.521044e-14, 3.535872e-14, 3.551697e-14, 3.552038e-14, 
    3.557119e-14, 3.57145e-14, 3.546826e-14, 3.623324e-14, 3.575987e-14, 
    3.505871e-14, 3.520216e-14, 3.52227e-14, 3.516708e-14, 3.554537e-14, 
    3.540808e-14, 3.577841e-14, 3.567815e-14, 3.584249e-14, 3.576078e-14, 
    3.574876e-14, 3.564396e-14, 3.557877e-14, 3.541435e-14, 3.528081e-14, 
    3.517511e-14, 3.519967e-14, 3.531583e-14, 3.552667e-14, 3.572667e-14, 
    3.568281e-14, 3.582995e-14, 3.544113e-14, 3.560392e-14, 3.554094e-14, 
    3.570524e-14, 3.534578e-14, 3.565174e-14, 3.526775e-14, 3.530134e-14, 
    3.540535e-14, 3.561499e-14, 3.566149e-14, 3.571111e-14, 3.568048e-14, 
    3.553205e-14, 3.550777e-14, 3.540281e-14, 3.537384e-14, 3.5294e-14, 
    3.522794e-14, 3.528828e-14, 3.535169e-14, 3.55321e-14, 3.569503e-14, 
    3.587306e-14, 3.59167e-14, 3.612527e-14, 3.59554e-14, 3.623587e-14, 
    3.59973e-14, 3.641077e-14, 3.566954e-14, 3.59904e-14, 3.54101e-14, 
    3.547241e-14, 3.558522e-14, 3.584463e-14, 3.57045e-14, 3.586842e-14, 
    3.550682e-14, 3.531984e-14, 3.527156e-14, 3.518153e-14, 3.527361e-14, 
    3.526612e-14, 3.535434e-14, 3.532597e-14, 3.553809e-14, 3.542408e-14, 
    3.574841e-14, 3.58671e-14, 3.620328e-14, 3.641006e-14, 3.662115e-14, 
    3.671451e-14, 3.674294e-14, 3.675483e-14 ;

 F_NIT =
  5.750217e-11, 5.781313e-11, 5.775263e-11, 5.800385e-11, 5.786444e-11, 
    5.802901e-11, 5.756515e-11, 5.782544e-11, 5.765922e-11, 5.753012e-11, 
    5.849272e-11, 5.801504e-11, 5.899102e-11, 5.868493e-11, 5.945526e-11, 
    5.894332e-11, 5.955875e-11, 5.944051e-11, 5.979681e-11, 5.969462e-11, 
    6.015131e-11, 5.984398e-11, 6.038875e-11, 6.007787e-11, 6.012642e-11, 
    5.983382e-11, 5.811111e-11, 5.843317e-11, 5.809203e-11, 5.81379e-11, 
    5.811732e-11, 5.786728e-11, 5.774143e-11, 5.747842e-11, 5.752613e-11, 
    5.771934e-11, 5.81585e-11, 5.800927e-11, 5.838576e-11, 5.837725e-11, 
    5.879765e-11, 5.860792e-11, 5.931663e-11, 5.911481e-11, 5.969888e-11, 
    5.955173e-11, 5.969195e-11, 5.964942e-11, 5.969249e-11, 5.947676e-11, 
    5.956913e-11, 5.937948e-11, 5.864348e-11, 5.885935e-11, 5.821654e-11, 
    5.783151e-11, 5.757652e-11, 5.739587e-11, 5.742138e-11, 5.747004e-11, 
    5.772046e-11, 5.795639e-11, 5.813648e-11, 5.825707e-11, 5.837602e-11, 
    5.873661e-11, 5.892799e-11, 5.935744e-11, 5.927987e-11, 5.941133e-11, 
    5.95371e-11, 5.974848e-11, 5.971366e-11, 5.980686e-11, 5.940787e-11, 
    5.967288e-11, 5.923566e-11, 5.935508e-11, 5.840826e-11, 5.804954e-11, 
    5.789725e-11, 5.77642e-11, 5.7441e-11, 5.766409e-11, 5.757609e-11, 
    5.778556e-11, 5.791883e-11, 5.78529e-11, 5.826037e-11, 5.810179e-11, 
    5.893933e-11, 5.85779e-11, 5.952243e-11, 5.929578e-11, 5.95768e-11, 
    5.943333e-11, 5.967924e-11, 5.94579e-11, 5.984158e-11, 5.992525e-11, 
    5.986805e-11, 6.008793e-11, 5.944561e-11, 5.969188e-11, 5.785108e-11, 
    5.786183e-11, 5.791192e-11, 5.769182e-11, 5.767837e-11, 5.747708e-11, 
    5.765617e-11, 5.773251e-11, 5.792656e-11, 5.804145e-11, 5.815077e-11, 
    5.839148e-11, 5.866082e-11, 5.903844e-11, 5.931045e-11, 5.949308e-11, 
    5.938107e-11, 5.947995e-11, 5.936941e-11, 5.931762e-11, 5.989387e-11, 
    5.956997e-11, 6.005627e-11, 6.002932e-11, 5.980904e-11, 6.003234e-11, 
    5.786937e-11, 5.780751e-11, 5.759297e-11, 5.776083e-11, 5.745516e-11, 
    5.762614e-11, 5.772455e-11, 5.810506e-11, 5.818885e-11, 5.826654e-11, 
    5.842018e-11, 5.861759e-11, 5.896465e-11, 5.926738e-11, 5.954441e-11, 
    5.952409e-11, 5.953123e-11, 5.959317e-11, 5.943977e-11, 5.961836e-11, 
    5.964834e-11, 5.956993e-11, 6.00257e-11, 5.989533e-11, 6.002873e-11, 
    5.994383e-11, 5.782761e-11, 5.793171e-11, 5.787544e-11, 5.798126e-11, 
    5.790668e-11, 5.823857e-11, 5.833824e-11, 5.880572e-11, 5.86137e-11, 
    5.891949e-11, 5.864472e-11, 5.869336e-11, 5.89294e-11, 5.865956e-11, 
    5.925063e-11, 5.884954e-11, 5.959556e-11, 5.919391e-11, 5.962077e-11, 
    5.954317e-11, 5.967168e-11, 5.978686e-11, 5.993194e-11, 6.020002e-11, 
    6.013789e-11, 6.036242e-11, 5.808708e-11, 5.822239e-11, 5.821049e-11, 
    5.835225e-11, 5.845719e-11, 5.868497e-11, 5.905113e-11, 5.891332e-11, 
    5.916644e-11, 5.92173e-11, 5.883279e-11, 5.906871e-11, 5.8313e-11, 
    5.843476e-11, 5.836226e-11, 5.809767e-11, 5.894497e-11, 5.850941e-11, 
    5.931489e-11, 5.907807e-11, 5.977041e-11, 5.94256e-11, 6.01037e-11, 
    6.039458e-11, 6.066907e-11, 6.099039e-11, 5.829632e-11, 5.82043e-11, 
    5.836913e-11, 5.859747e-11, 5.880978e-11, 5.909255e-11, 5.912153e-11, 
    5.917457e-11, 5.93121e-11, 5.942784e-11, 5.91913e-11, 5.945686e-11, 
    5.846295e-11, 5.898286e-11, 5.816944e-11, 5.841379e-11, 5.858394e-11, 
    5.85093e-11, 5.889752e-11, 5.898917e-11, 5.93623e-11, 5.916929e-11, 
    6.032268e-11, 5.981113e-11, 6.123567e-11, 6.083601e-11, 5.817216e-11, 
    5.8296e-11, 5.872794e-11, 5.852224e-11, 5.911145e-11, 5.925688e-11, 
    5.937525e-11, 5.952668e-11, 5.954305e-11, 5.963287e-11, 5.94857e-11, 
    5.962705e-11, 5.90931e-11, 5.933144e-11, 5.867847e-11, 5.883707e-11, 
    5.876409e-11, 5.868406e-11, 5.893119e-11, 5.919495e-11, 5.920064e-11, 
    5.928532e-11, 5.952417e-11, 5.911376e-11, 6.038874e-11, 5.959979e-11, 
    5.843118e-11, 5.867026e-11, 5.87045e-11, 5.86118e-11, 5.924228e-11, 
    5.901347e-11, 5.963068e-11, 5.946359e-11, 5.973748e-11, 5.96013e-11, 
    5.958126e-11, 5.94066e-11, 5.929796e-11, 5.902391e-11, 5.880135e-11, 
    5.862519e-11, 5.866613e-11, 5.885972e-11, 5.921111e-11, 5.954445e-11, 
    5.947134e-11, 5.971658e-11, 5.906854e-11, 5.933986e-11, 5.92349e-11, 
    5.950873e-11, 5.890963e-11, 5.941956e-11, 5.877958e-11, 5.883557e-11, 
    5.900892e-11, 5.935832e-11, 5.943581e-11, 5.951852e-11, 5.946747e-11, 
    5.922009e-11, 5.917961e-11, 5.900468e-11, 5.89564e-11, 5.882334e-11, 
    5.871324e-11, 5.881381e-11, 5.891948e-11, 5.922017e-11, 5.949172e-11, 
    5.978843e-11, 5.986117e-11, 6.020878e-11, 5.992568e-11, 6.039312e-11, 
    5.999549e-11, 6.068461e-11, 5.944924e-11, 5.9984e-11, 5.901683e-11, 
    5.912069e-11, 5.93087e-11, 5.974105e-11, 5.95075e-11, 5.978069e-11, 
    5.917803e-11, 5.886639e-11, 5.878593e-11, 5.863588e-11, 5.878936e-11, 
    5.877687e-11, 5.892389e-11, 5.887662e-11, 5.923016e-11, 5.904013e-11, 
    5.958068e-11, 5.977849e-11, 6.03388e-11, 6.068343e-11, 6.103525e-11, 
    6.119084e-11, 6.123824e-11, 6.125805e-11 ;

 F_NIT_vr =
  2.588892e-10, 2.599761e-10, 2.597642e-10, 2.606412e-10, 2.601545e-10, 
    2.607282e-10, 2.591083e-10, 2.600172e-10, 2.594366e-10, 2.589849e-10, 
    2.623419e-10, 2.606782e-10, 2.64074e-10, 2.630105e-10, 2.656828e-10, 
    2.639076e-10, 2.660408e-10, 2.656313e-10, 2.668639e-10, 2.665103e-10, 
    2.680869e-10, 2.670263e-10, 2.689052e-10, 2.678333e-10, 2.680003e-10, 
    2.669899e-10, 2.610152e-10, 2.621366e-10, 2.609482e-10, 2.611081e-10, 
    2.610361e-10, 2.601632e-10, 2.597234e-10, 2.588039e-10, 2.589704e-10, 
    2.596457e-10, 2.61178e-10, 2.606574e-10, 2.619693e-10, 2.619397e-10, 
    2.634013e-10, 2.627419e-10, 2.652019e-10, 2.645018e-10, 2.665247e-10, 
    2.660152e-10, 2.665002e-10, 2.663527e-10, 2.665013e-10, 2.657548e-10, 
    2.660739e-10, 2.654174e-10, 2.628686e-10, 2.636184e-10, 2.613817e-10, 
    2.600377e-10, 2.591469e-10, 2.585151e-10, 2.586038e-10, 2.58774e-10, 
    2.596491e-10, 2.604727e-10, 2.611008e-10, 2.615207e-10, 2.619346e-10, 
    2.631885e-10, 2.638533e-10, 2.653425e-10, 2.650738e-10, 2.655287e-10, 
    2.659642e-10, 2.66695e-10, 2.665746e-10, 2.668963e-10, 2.655155e-10, 
    2.664327e-10, 2.649183e-10, 2.653322e-10, 2.620485e-10, 2.60799e-10, 
    2.60267e-10, 2.598024e-10, 2.586722e-10, 2.594523e-10, 2.591443e-10, 
    2.598761e-10, 2.603413e-10, 2.601108e-10, 2.615319e-10, 2.609787e-10, 
    2.638923e-10, 2.626364e-10, 2.659138e-10, 2.651284e-10, 2.661013e-10, 
    2.656047e-10, 2.66455e-10, 2.656892e-10, 2.670157e-10, 2.673048e-10, 
    2.671066e-10, 2.678661e-10, 2.65645e-10, 2.664972e-10, 2.601059e-10, 
    2.601435e-10, 2.60318e-10, 2.595487e-10, 2.595017e-10, 2.587976e-10, 
    2.594235e-10, 2.596902e-10, 2.603676e-10, 2.60768e-10, 2.611489e-10, 
    2.619876e-10, 2.629242e-10, 2.642356e-10, 2.651789e-10, 2.658112e-10, 
    2.654232e-10, 2.657652e-10, 2.653822e-10, 2.652024e-10, 2.671955e-10, 
    2.660757e-10, 2.67756e-10, 2.676631e-10, 2.669017e-10, 2.676727e-10, 
    2.601693e-10, 2.599529e-10, 2.592031e-10, 2.597894e-10, 2.587204e-10, 
    2.593183e-10, 2.596617e-10, 2.609895e-10, 2.612815e-10, 2.615522e-10, 
    2.62087e-10, 2.627735e-10, 2.639792e-10, 2.65029e-10, 2.659885e-10, 
    2.659178e-10, 2.659424e-10, 2.661562e-10, 2.656251e-10, 2.662429e-10, 
    2.663462e-10, 2.660751e-10, 2.676498e-10, 2.671997e-10, 2.6766e-10, 
    2.673664e-10, 2.600228e-10, 2.603858e-10, 2.60189e-10, 2.605584e-10, 
    2.602975e-10, 2.614549e-10, 2.618017e-10, 2.634275e-10, 2.627599e-10, 
    2.638225e-10, 2.628673e-10, 2.630364e-10, 2.638556e-10, 2.629183e-10, 
    2.649699e-10, 2.635775e-10, 2.661643e-10, 2.64772e-10, 2.662509e-10, 
    2.659821e-10, 2.664263e-10, 2.668246e-10, 2.673253e-10, 2.682504e-10, 
    2.680356e-10, 2.688099e-10, 2.609276e-10, 2.613987e-10, 2.613574e-10, 
    2.618508e-10, 2.622157e-10, 2.630082e-10, 2.642795e-10, 2.638009e-10, 
    2.646789e-10, 2.648553e-10, 2.635204e-10, 2.643393e-10, 2.617117e-10, 
    2.621351e-10, 2.618829e-10, 2.609603e-10, 2.639083e-10, 2.623939e-10, 
    2.651911e-10, 2.643696e-10, 2.667669e-10, 2.655737e-10, 2.679175e-10, 
    2.689201e-10, 2.698652e-10, 2.709688e-10, 2.616561e-10, 2.613352e-10, 
    2.619091e-10, 2.627035e-10, 2.634412e-10, 2.644229e-10, 2.645232e-10, 
    2.647067e-10, 2.651832e-10, 2.655842e-10, 2.647639e-10, 2.656839e-10, 
    2.622325e-10, 2.640399e-10, 2.612101e-10, 2.620611e-10, 2.626528e-10, 
    2.623933e-10, 2.637427e-10, 2.640605e-10, 2.653538e-10, 2.646851e-10, 
    2.686715e-10, 2.669062e-10, 2.718104e-10, 2.704381e-10, 2.612228e-10, 
    2.61654e-10, 2.631564e-10, 2.624413e-10, 2.644878e-10, 2.649921e-10, 
    2.654018e-10, 2.659261e-10, 2.659823e-10, 2.66293e-10, 2.657833e-10, 
    2.662725e-10, 2.64422e-10, 2.652485e-10, 2.629819e-10, 2.635325e-10, 
    2.63279e-10, 2.630004e-10, 2.638587e-10, 2.647736e-10, 2.647932e-10, 
    2.650862e-10, 2.659123e-10, 2.64491e-10, 2.688975e-10, 2.661733e-10, 
    2.621245e-10, 2.629554e-10, 2.630744e-10, 2.627522e-10, 2.649408e-10, 
    2.641471e-10, 2.662855e-10, 2.657068e-10, 2.666542e-10, 2.661832e-10, 
    2.661133e-10, 2.655087e-10, 2.651317e-10, 2.641812e-10, 2.634079e-10, 
    2.627957e-10, 2.629375e-10, 2.636102e-10, 2.648289e-10, 2.659838e-10, 
    2.657303e-10, 2.665786e-10, 2.643336e-10, 2.652742e-10, 2.649098e-10, 
    2.658587e-10, 2.637869e-10, 2.655545e-10, 2.63335e-10, 2.635291e-10, 
    2.641306e-10, 2.653419e-10, 2.656101e-10, 2.658964e-10, 2.657193e-10, 
    2.64862e-10, 2.647214e-10, 2.641143e-10, 2.639462e-10, 2.634843e-10, 
    2.631011e-10, 2.634506e-10, 2.638169e-10, 2.648604e-10, 2.658007e-10, 
    2.668267e-10, 2.670781e-10, 2.682769e-10, 2.672998e-10, 2.689112e-10, 
    2.675396e-10, 2.699146e-10, 2.656569e-10, 2.67506e-10, 2.641582e-10, 
    2.645181e-10, 2.651695e-10, 2.666656e-10, 2.658576e-10, 2.668024e-10, 
    2.647158e-10, 2.636336e-10, 2.63354e-10, 2.628325e-10, 2.633654e-10, 
    2.633221e-10, 2.638325e-10, 2.636679e-10, 2.648942e-10, 2.642353e-10, 
    2.661077e-10, 2.667918e-10, 2.687253e-10, 2.699114e-10, 2.711207e-10, 
    2.716543e-10, 2.718168e-10, 2.718844e-10,
  1.737267e-10, 1.746417e-10, 1.744638e-10, 1.752024e-10, 1.747927e-10, 
    1.752764e-10, 1.739122e-10, 1.746779e-10, 1.741891e-10, 1.738092e-10, 
    1.766379e-10, 1.752354e-10, 1.780994e-10, 1.772023e-10, 1.794585e-10, 
    1.779595e-10, 1.797613e-10, 1.794156e-10, 1.804574e-10, 1.801588e-10, 
    1.814923e-10, 1.805953e-10, 1.821852e-10, 1.812782e-10, 1.814199e-10, 
    1.805656e-10, 1.755177e-10, 1.76463e-10, 1.754617e-10, 1.755964e-10, 
    1.75536e-10, 1.74801e-10, 1.744308e-10, 1.73657e-10, 1.737975e-10, 
    1.743659e-10, 1.75657e-10, 1.752187e-10, 1.763246e-10, 1.762996e-10, 
    1.775329e-10, 1.769765e-10, 1.790531e-10, 1.784624e-10, 1.801713e-10, 
    1.79741e-10, 1.80151e-10, 1.800267e-10, 1.801526e-10, 1.795218e-10, 
    1.79792e-10, 1.792372e-10, 1.770806e-10, 1.777136e-10, 1.758275e-10, 
    1.746956e-10, 1.739457e-10, 1.734139e-10, 1.734891e-10, 1.736323e-10, 
    1.743693e-10, 1.750632e-10, 1.755925e-10, 1.759468e-10, 1.76296e-10, 
    1.773536e-10, 1.779148e-10, 1.791725e-10, 1.789456e-10, 1.793302e-10, 
    1.796983e-10, 1.803162e-10, 1.802145e-10, 1.804868e-10, 1.793203e-10, 
    1.800953e-10, 1.788164e-10, 1.791659e-10, 1.763899e-10, 1.753369e-10, 
    1.74889e-10, 1.744979e-10, 1.735469e-10, 1.742034e-10, 1.739445e-10, 
    1.745609e-10, 1.749528e-10, 1.74759e-10, 1.759564e-10, 1.754906e-10, 
    1.779481e-10, 1.768884e-10, 1.796553e-10, 1.789922e-10, 1.798144e-10, 
    1.793948e-10, 1.801138e-10, 1.794667e-10, 1.805883e-10, 1.808327e-10, 
    1.806656e-10, 1.813078e-10, 1.794308e-10, 1.801509e-10, 1.747535e-10, 
    1.747851e-10, 1.749325e-10, 1.74285e-10, 1.742455e-10, 1.736531e-10, 
    1.741803e-10, 1.744048e-10, 1.749756e-10, 1.753133e-10, 1.756345e-10, 
    1.763414e-10, 1.771316e-10, 1.782386e-10, 1.790352e-10, 1.795696e-10, 
    1.792419e-10, 1.795312e-10, 1.792078e-10, 1.790563e-10, 1.80741e-10, 
    1.797944e-10, 1.812154e-10, 1.811368e-10, 1.804933e-10, 1.811456e-10, 
    1.748073e-10, 1.746255e-10, 1.739942e-10, 1.744882e-10, 1.735887e-10, 
    1.740919e-10, 1.743813e-10, 1.755001e-10, 1.757464e-10, 1.759746e-10, 
    1.764257e-10, 1.77005e-10, 1.780224e-10, 1.789091e-10, 1.797197e-10, 
    1.796603e-10, 1.796812e-10, 1.798623e-10, 1.794137e-10, 1.79936e-10, 
    1.800236e-10, 1.797944e-10, 1.811262e-10, 1.807455e-10, 1.811351e-10, 
    1.808872e-10, 1.746846e-10, 1.749907e-10, 1.748253e-10, 1.751363e-10, 
    1.749171e-10, 1.758923e-10, 1.761849e-10, 1.775565e-10, 1.769935e-10, 
    1.7789e-10, 1.770846e-10, 1.772272e-10, 1.779188e-10, 1.771282e-10, 
    1.7886e-10, 1.77685e-10, 1.798694e-10, 1.786938e-10, 1.799431e-10, 
    1.797162e-10, 1.80092e-10, 1.804286e-10, 1.808524e-10, 1.816349e-10, 
    1.814537e-10, 1.821088e-10, 1.754474e-10, 1.758448e-10, 1.7581e-10, 
    1.762263e-10, 1.765343e-10, 1.772027e-10, 1.782758e-10, 1.778721e-10, 
    1.786137e-10, 1.787626e-10, 1.776362e-10, 1.783273e-10, 1.761111e-10, 
    1.764684e-10, 1.762558e-10, 1.754786e-10, 1.779648e-10, 1.766876e-10, 
    1.790483e-10, 1.78355e-10, 1.803805e-10, 1.793722e-10, 1.813539e-10, 
    1.822022e-10, 1.830026e-10, 1.839379e-10, 1.76062e-10, 1.757919e-10, 
    1.762759e-10, 1.769458e-10, 1.775686e-10, 1.783972e-10, 1.784821e-10, 
    1.786374e-10, 1.790401e-10, 1.793788e-10, 1.786863e-10, 1.794637e-10, 
    1.765509e-10, 1.780759e-10, 1.756896e-10, 1.764069e-10, 1.769064e-10, 
    1.766875e-10, 1.778261e-10, 1.780947e-10, 1.791871e-10, 1.786223e-10, 
    1.819926e-10, 1.804994e-10, 1.846515e-10, 1.834886e-10, 1.756974e-10, 
    1.760612e-10, 1.773286e-10, 1.767253e-10, 1.784527e-10, 1.788784e-10, 
    1.79225e-10, 1.796678e-10, 1.797158e-10, 1.799784e-10, 1.795481e-10, 
    1.799615e-10, 1.783989e-10, 1.790968e-10, 1.771838e-10, 1.776488e-10, 
    1.774349e-10, 1.772003e-10, 1.779248e-10, 1.786972e-10, 1.78714e-10, 
    1.789618e-10, 1.7966e-10, 1.784597e-10, 1.821848e-10, 1.798813e-10, 
    1.764581e-10, 1.771593e-10, 1.7726e-10, 1.769881e-10, 1.788357e-10, 
    1.781656e-10, 1.799721e-10, 1.794834e-10, 1.802843e-10, 1.798862e-10, 
    1.798276e-10, 1.793168e-10, 1.789988e-10, 1.781963e-10, 1.775441e-10, 
    1.770276e-10, 1.771477e-10, 1.777152e-10, 1.787445e-10, 1.7972e-10, 
    1.795062e-10, 1.802234e-10, 1.783272e-10, 1.791215e-10, 1.788143e-10, 
    1.796157e-10, 1.778614e-10, 1.793539e-10, 1.774802e-10, 1.776444e-10, 
    1.781524e-10, 1.791752e-10, 1.794022e-10, 1.79644e-10, 1.794949e-10, 
    1.787707e-10, 1.786523e-10, 1.781401e-10, 1.779985e-10, 1.776087e-10, 
    1.772859e-10, 1.775807e-10, 1.778904e-10, 1.787712e-10, 1.795658e-10, 
    1.804333e-10, 1.806459e-10, 1.816603e-10, 1.808339e-10, 1.821976e-10, 
    1.810373e-10, 1.830475e-10, 1.79441e-10, 1.810039e-10, 1.781756e-10, 
    1.784798e-10, 1.7903e-10, 1.802945e-10, 1.796119e-10, 1.804104e-10, 
    1.786477e-10, 1.777346e-10, 1.77499e-10, 1.770589e-10, 1.775091e-10, 
    1.774725e-10, 1.779035e-10, 1.77765e-10, 1.788005e-10, 1.78244e-10, 
    1.798261e-10, 1.804042e-10, 1.8204e-10, 1.830444e-10, 1.840688e-10, 
    1.845214e-10, 1.846592e-10, 1.847168e-10,
  1.861625e-10, 1.871557e-10, 1.869625e-10, 1.877644e-10, 1.873196e-10, 
    1.878448e-10, 1.863638e-10, 1.87195e-10, 1.866643e-10, 1.86252e-10, 
    1.893236e-10, 1.878003e-10, 1.909113e-10, 1.899365e-10, 1.923887e-10, 
    1.907594e-10, 1.927178e-10, 1.923419e-10, 1.934747e-10, 1.9315e-10, 
    1.946005e-10, 1.936246e-10, 1.953542e-10, 1.943675e-10, 1.945216e-10, 
    1.935924e-10, 1.881068e-10, 1.891336e-10, 1.880459e-10, 1.881923e-10, 
    1.881266e-10, 1.873287e-10, 1.869267e-10, 1.860868e-10, 1.862393e-10, 
    1.868563e-10, 1.882581e-10, 1.87782e-10, 1.889831e-10, 1.889559e-10, 
    1.902957e-10, 1.896912e-10, 1.919479e-10, 1.913057e-10, 1.931635e-10, 
    1.926957e-10, 1.931415e-10, 1.930063e-10, 1.931432e-10, 1.924573e-10, 
    1.927511e-10, 1.92148e-10, 1.898043e-10, 1.904921e-10, 1.884432e-10, 
    1.872143e-10, 1.864002e-10, 1.85823e-10, 1.859046e-10, 1.8606e-10, 
    1.868599e-10, 1.876133e-10, 1.88188e-10, 1.885727e-10, 1.88952e-10, 
    1.90101e-10, 1.907107e-10, 1.920777e-10, 1.91831e-10, 1.922491e-10, 
    1.926492e-10, 1.933212e-10, 1.932105e-10, 1.935067e-10, 1.922383e-10, 
    1.930809e-10, 1.916905e-10, 1.920704e-10, 1.890542e-10, 1.879105e-10, 
    1.874242e-10, 1.869996e-10, 1.859673e-10, 1.866799e-10, 1.863989e-10, 
    1.870679e-10, 1.874934e-10, 1.87283e-10, 1.885832e-10, 1.880773e-10, 
    1.907469e-10, 1.895955e-10, 1.926025e-10, 1.918816e-10, 1.927755e-10, 
    1.923193e-10, 1.931011e-10, 1.923974e-10, 1.936171e-10, 1.938829e-10, 
    1.937012e-10, 1.943996e-10, 1.923584e-10, 1.931414e-10, 1.87277e-10, 
    1.873113e-10, 1.874713e-10, 1.867685e-10, 1.867256e-10, 1.860826e-10, 
    1.866547e-10, 1.868985e-10, 1.875181e-10, 1.878848e-10, 1.882336e-10, 
    1.890013e-10, 1.898598e-10, 1.910626e-10, 1.919283e-10, 1.925093e-10, 
    1.921531e-10, 1.924676e-10, 1.92116e-10, 1.919513e-10, 1.937832e-10, 
    1.927538e-10, 1.942991e-10, 1.942136e-10, 1.935137e-10, 1.942232e-10, 
    1.873354e-10, 1.87138e-10, 1.864528e-10, 1.86989e-10, 1.860126e-10, 
    1.865588e-10, 1.868731e-10, 1.880877e-10, 1.883551e-10, 1.886029e-10, 
    1.890929e-10, 1.897221e-10, 1.908276e-10, 1.917913e-10, 1.926725e-10, 
    1.926079e-10, 1.926307e-10, 1.928276e-10, 1.923398e-10, 1.929077e-10, 
    1.93003e-10, 1.927538e-10, 1.942021e-10, 1.93788e-10, 1.942117e-10, 
    1.939421e-10, 1.872022e-10, 1.875345e-10, 1.873549e-10, 1.876927e-10, 
    1.874546e-10, 1.885136e-10, 1.888315e-10, 1.903214e-10, 1.897097e-10, 
    1.906838e-10, 1.898086e-10, 1.899636e-10, 1.907152e-10, 1.89856e-10, 
    1.917379e-10, 1.90461e-10, 1.928352e-10, 1.915574e-10, 1.929154e-10, 
    1.926687e-10, 1.930773e-10, 1.934433e-10, 1.939043e-10, 1.947555e-10, 
    1.945584e-10, 1.952711e-10, 1.880304e-10, 1.88462e-10, 1.884242e-10, 
    1.888763e-10, 1.892108e-10, 1.899369e-10, 1.91103e-10, 1.906643e-10, 
    1.914701e-10, 1.91632e-10, 1.904079e-10, 1.91159e-10, 1.887512e-10, 
    1.891393e-10, 1.889083e-10, 1.880643e-10, 1.907651e-10, 1.893774e-10, 
    1.919426e-10, 1.91189e-10, 1.933911e-10, 1.922948e-10, 1.944498e-10, 
    1.953729e-10, 1.962438e-10, 1.97262e-10, 1.886979e-10, 1.884044e-10, 
    1.889301e-10, 1.896579e-10, 1.903345e-10, 1.912349e-10, 1.913272e-10, 
    1.91496e-10, 1.919337e-10, 1.923019e-10, 1.915492e-10, 1.923942e-10, 
    1.892291e-10, 1.908858e-10, 1.882934e-10, 1.890725e-10, 1.896151e-10, 
    1.893772e-10, 1.906142e-10, 1.909061e-10, 1.920935e-10, 1.914795e-10, 
    1.951448e-10, 1.935204e-10, 1.98039e-10, 1.967729e-10, 1.883019e-10, 
    1.88697e-10, 1.900737e-10, 1.894183e-10, 1.912951e-10, 1.91758e-10, 
    1.921346e-10, 1.926161e-10, 1.926683e-10, 1.929538e-10, 1.92486e-10, 
    1.929354e-10, 1.912368e-10, 1.919953e-10, 1.899164e-10, 1.904216e-10, 
    1.901892e-10, 1.899342e-10, 1.907215e-10, 1.91561e-10, 1.915792e-10, 
    1.918486e-10, 1.926079e-10, 1.913028e-10, 1.953542e-10, 1.928485e-10, 
    1.89128e-10, 1.898899e-10, 1.899991e-10, 1.897038e-10, 1.917115e-10, 
    1.909832e-10, 1.929469e-10, 1.924156e-10, 1.932864e-10, 1.928535e-10, 
    1.927898e-10, 1.922344e-10, 1.918888e-10, 1.910166e-10, 1.903079e-10, 
    1.897467e-10, 1.898771e-10, 1.904938e-10, 1.916125e-10, 1.926729e-10, 
    1.924404e-10, 1.932202e-10, 1.911589e-10, 1.920222e-10, 1.916883e-10, 
    1.925594e-10, 1.906526e-10, 1.922751e-10, 1.902384e-10, 1.904168e-10, 
    1.909688e-10, 1.920806e-10, 1.923273e-10, 1.925903e-10, 1.92428e-10, 
    1.91641e-10, 1.915122e-10, 1.909554e-10, 1.908017e-10, 1.90378e-10, 
    1.900273e-10, 1.903476e-10, 1.906841e-10, 1.916414e-10, 1.925052e-10, 
    1.934485e-10, 1.936797e-10, 1.947833e-10, 1.938844e-10, 1.953681e-10, 
    1.941058e-10, 1.962929e-10, 1.923697e-10, 1.940693e-10, 1.90994e-10, 
    1.913247e-10, 1.919228e-10, 1.932976e-10, 1.925553e-10, 1.934237e-10, 
    1.915072e-10, 1.90515e-10, 1.902588e-10, 1.897807e-10, 1.902697e-10, 
    1.9023e-10, 1.906983e-10, 1.905478e-10, 1.916732e-10, 1.910684e-10, 
    1.927882e-10, 1.934169e-10, 1.951962e-10, 1.962893e-10, 1.974045e-10, 
    1.978973e-10, 1.980474e-10, 1.981101e-10,
  1.982555e-10, 1.993355e-10, 1.991255e-10, 1.999979e-10, 1.995138e-10, 
    2.000853e-10, 1.984744e-10, 1.993784e-10, 1.988011e-10, 1.983528e-10, 
    2.016953e-10, 2.000369e-10, 2.034247e-10, 2.023625e-10, 2.050355e-10, 
    2.032592e-10, 2.053945e-10, 2.049844e-10, 2.062202e-10, 2.058659e-10, 
    2.074496e-10, 2.063839e-10, 2.082728e-10, 2.07195e-10, 2.073633e-10, 
    2.063487e-10, 2.003703e-10, 2.014885e-10, 2.003041e-10, 2.004634e-10, 
    2.003919e-10, 1.995237e-10, 1.990867e-10, 1.981732e-10, 1.983389e-10, 
    1.9901e-10, 2.00535e-10, 2.000169e-10, 2.013241e-10, 2.012946e-10, 
    2.027538e-10, 2.020953e-10, 2.045546e-10, 2.038544e-10, 2.058806e-10, 
    2.053703e-10, 2.058567e-10, 2.057091e-10, 2.058586e-10, 2.051103e-10, 
    2.054307e-10, 2.047728e-10, 2.022185e-10, 2.029678e-10, 2.007364e-10, 
    1.993995e-10, 1.985139e-10, 1.978864e-10, 1.979751e-10, 1.981441e-10, 
    1.990139e-10, 1.998333e-10, 2.004586e-10, 2.008773e-10, 2.012903e-10, 
    2.02542e-10, 2.032062e-10, 2.046962e-10, 2.044272e-10, 2.048832e-10, 
    2.053196e-10, 2.060527e-10, 2.05932e-10, 2.062552e-10, 2.048713e-10, 
    2.057906e-10, 2.042739e-10, 2.046883e-10, 2.01402e-10, 2.001567e-10, 
    1.996278e-10, 1.991658e-10, 1.980433e-10, 1.988181e-10, 1.985125e-10, 
    1.992401e-10, 1.997029e-10, 1.99474e-10, 2.008888e-10, 2.003382e-10, 
    2.032455e-10, 2.019911e-10, 2.052686e-10, 2.044824e-10, 2.054573e-10, 
    2.049596e-10, 2.058126e-10, 2.050449e-10, 2.063757e-10, 2.066659e-10, 
    2.064675e-10, 2.0723e-10, 2.050023e-10, 2.058566e-10, 1.994675e-10, 
    1.995048e-10, 1.996788e-10, 1.989145e-10, 1.988678e-10, 1.981686e-10, 
    1.987907e-10, 1.990559e-10, 1.997298e-10, 2.001287e-10, 2.005084e-10, 
    2.01344e-10, 2.02279e-10, 2.035895e-10, 2.045333e-10, 2.051669e-10, 
    2.047783e-10, 2.051214e-10, 2.047379e-10, 2.045583e-10, 2.06557e-10, 
    2.054337e-10, 2.071203e-10, 2.070268e-10, 2.062629e-10, 2.070373e-10, 
    1.995311e-10, 1.993163e-10, 1.985712e-10, 1.991542e-10, 1.980926e-10, 
    1.986864e-10, 1.990282e-10, 2.003496e-10, 2.006406e-10, 2.009103e-10, 
    2.014437e-10, 2.02129e-10, 2.033335e-10, 2.043839e-10, 2.05345e-10, 
    2.052745e-10, 2.052993e-10, 2.055142e-10, 2.04982e-10, 2.056016e-10, 
    2.057056e-10, 2.054336e-10, 2.070143e-10, 2.065622e-10, 2.070248e-10, 
    2.067305e-10, 1.993861e-10, 1.997476e-10, 1.995522e-10, 1.999197e-10, 
    1.996608e-10, 2.008131e-10, 2.011592e-10, 2.027819e-10, 2.021154e-10, 
    2.031767e-10, 2.022232e-10, 2.02392e-10, 2.032112e-10, 2.022747e-10, 
    2.043258e-10, 2.029341e-10, 2.055225e-10, 2.041291e-10, 2.056099e-10, 
    2.053408e-10, 2.057866e-10, 2.061861e-10, 2.066892e-10, 2.076187e-10, 
    2.074034e-10, 2.081818e-10, 2.002872e-10, 2.00757e-10, 2.007157e-10, 
    2.012079e-10, 2.015722e-10, 2.023628e-10, 2.036335e-10, 2.031554e-10, 
    2.040337e-10, 2.042102e-10, 2.02876e-10, 2.036946e-10, 2.010717e-10, 
    2.014944e-10, 2.012428e-10, 2.003242e-10, 2.032653e-10, 2.017536e-10, 
    2.045489e-10, 2.037273e-10, 2.061291e-10, 2.04933e-10, 2.072848e-10, 
    2.082933e-10, 2.092448e-10, 2.103583e-10, 2.010137e-10, 2.006942e-10, 
    2.012665e-10, 2.020591e-10, 2.027961e-10, 2.037773e-10, 2.038779e-10, 
    2.040619e-10, 2.045391e-10, 2.049406e-10, 2.0412e-10, 2.050413e-10, 
    2.015923e-10, 2.033968e-10, 2.005734e-10, 2.014217e-10, 2.020124e-10, 
    2.017533e-10, 2.031008e-10, 2.034189e-10, 2.047135e-10, 2.040439e-10, 
    2.080441e-10, 2.062703e-10, 2.112082e-10, 2.098234e-10, 2.005826e-10, 
    2.010126e-10, 2.02512e-10, 2.017981e-10, 2.038429e-10, 2.043475e-10, 
    2.047582e-10, 2.052835e-10, 2.053404e-10, 2.056519e-10, 2.051415e-10, 
    2.056317e-10, 2.037794e-10, 2.046063e-10, 2.023405e-10, 2.02891e-10, 
    2.026377e-10, 2.0236e-10, 2.032177e-10, 2.041329e-10, 2.041527e-10, 
    2.044465e-10, 2.05275e-10, 2.038513e-10, 2.082731e-10, 2.055374e-10, 
    2.01482e-10, 2.023118e-10, 2.024307e-10, 2.02109e-10, 2.042969e-10, 
    2.03503e-10, 2.056443e-10, 2.050647e-10, 2.060148e-10, 2.055424e-10, 
    2.05473e-10, 2.048671e-10, 2.044902e-10, 2.035394e-10, 2.027671e-10, 
    2.021556e-10, 2.022978e-10, 2.029697e-10, 2.04189e-10, 2.053454e-10, 
    2.050918e-10, 2.059425e-10, 2.036944e-10, 2.046357e-10, 2.042717e-10, 
    2.052216e-10, 2.031426e-10, 2.049119e-10, 2.026913e-10, 2.028857e-10, 
    2.034873e-10, 2.046995e-10, 2.049684e-10, 2.052553e-10, 2.050783e-10, 
    2.0422e-10, 2.040796e-10, 2.034727e-10, 2.033051e-10, 2.028434e-10, 
    2.024613e-10, 2.028103e-10, 2.031771e-10, 2.042204e-10, 2.051625e-10, 
    2.061917e-10, 2.06444e-10, 2.076493e-10, 2.066677e-10, 2.082884e-10, 
    2.069098e-10, 2.092988e-10, 2.050149e-10, 2.068696e-10, 2.035147e-10, 
    2.038751e-10, 2.045274e-10, 2.060272e-10, 2.052171e-10, 2.061647e-10, 
    2.040741e-10, 2.029928e-10, 2.027136e-10, 2.021928e-10, 2.027255e-10, 
    2.026821e-10, 2.031924e-10, 2.030284e-10, 2.042551e-10, 2.035958e-10, 
    2.054712e-10, 2.061573e-10, 2.081001e-10, 2.092947e-10, 2.10514e-10, 
    2.110531e-10, 2.112173e-10, 2.112859e-10,
  2.010477e-10, 2.02185e-10, 2.019636e-10, 2.02883e-10, 2.023727e-10, 
    2.029751e-10, 2.01278e-10, 2.022302e-10, 2.01622e-10, 2.011499e-10, 
    2.046739e-10, 2.029241e-10, 2.065008e-10, 2.053781e-10, 2.082051e-10, 
    2.063259e-10, 2.085852e-10, 2.081508e-10, 2.094601e-10, 2.090845e-10, 
    2.107643e-10, 2.096335e-10, 2.116381e-10, 2.104939e-10, 2.106726e-10, 
    2.095963e-10, 2.032755e-10, 2.044555e-10, 2.032057e-10, 2.033737e-10, 
    2.032983e-10, 2.023832e-10, 2.019229e-10, 2.009609e-10, 2.011354e-10, 
    2.01842e-10, 2.034493e-10, 2.029029e-10, 2.042816e-10, 2.042504e-10, 
    2.057914e-10, 2.050958e-10, 2.076959e-10, 2.06955e-10, 2.091002e-10, 
    2.085595e-10, 2.090748e-10, 2.089184e-10, 2.090768e-10, 2.082841e-10, 
    2.086235e-10, 2.079268e-10, 2.05226e-10, 2.060176e-10, 2.036617e-10, 
    2.022525e-10, 2.013197e-10, 2.006592e-10, 2.007525e-10, 2.009304e-10, 
    2.018462e-10, 2.027094e-10, 2.033686e-10, 2.038102e-10, 2.042459e-10, 
    2.055679e-10, 2.062697e-10, 2.078459e-10, 2.075609e-10, 2.080438e-10, 
    2.085057e-10, 2.092826e-10, 2.091546e-10, 2.094973e-10, 2.080311e-10, 
    2.090048e-10, 2.073987e-10, 2.078373e-10, 2.043644e-10, 2.030503e-10, 
    2.024931e-10, 2.020061e-10, 2.008243e-10, 2.0164e-10, 2.013182e-10, 
    2.020843e-10, 2.025719e-10, 2.023307e-10, 2.038223e-10, 2.032417e-10, 
    2.063113e-10, 2.049859e-10, 2.084518e-10, 2.076194e-10, 2.086516e-10, 
    2.081245e-10, 2.090281e-10, 2.082148e-10, 2.096249e-10, 2.099326e-10, 
    2.097223e-10, 2.10531e-10, 2.081698e-10, 2.090747e-10, 2.023239e-10, 
    2.023633e-10, 2.025466e-10, 2.017415e-10, 2.016922e-10, 2.009562e-10, 
    2.016111e-10, 2.018903e-10, 2.026002e-10, 2.030208e-10, 2.034211e-10, 
    2.043027e-10, 2.052899e-10, 2.066749e-10, 2.076733e-10, 2.083441e-10, 
    2.079326e-10, 2.082959e-10, 2.078898e-10, 2.076997e-10, 2.098173e-10, 
    2.086267e-10, 2.104146e-10, 2.103154e-10, 2.095054e-10, 2.103266e-10, 
    2.023909e-10, 2.021646e-10, 2.013799e-10, 2.019938e-10, 2.008761e-10, 
    2.015013e-10, 2.018613e-10, 2.032538e-10, 2.035605e-10, 2.038451e-10, 
    2.044078e-10, 2.051314e-10, 2.064042e-10, 2.075153e-10, 2.085326e-10, 
    2.08458e-10, 2.084843e-10, 2.087119e-10, 2.081483e-10, 2.088045e-10, 
    2.089147e-10, 2.086266e-10, 2.103021e-10, 2.098226e-10, 2.103133e-10, 
    2.10001e-10, 2.022381e-10, 2.026191e-10, 2.024132e-10, 2.028005e-10, 
    2.025276e-10, 2.037427e-10, 2.041078e-10, 2.058213e-10, 2.051171e-10, 
    2.062385e-10, 2.052309e-10, 2.054092e-10, 2.062751e-10, 2.052853e-10, 
    2.074539e-10, 2.059822e-10, 2.087207e-10, 2.072459e-10, 2.088134e-10, 
    2.085282e-10, 2.090004e-10, 2.094239e-10, 2.099573e-10, 2.109437e-10, 
    2.10715e-10, 2.115414e-10, 2.031878e-10, 2.036833e-10, 2.036397e-10, 
    2.04159e-10, 2.045435e-10, 2.053784e-10, 2.067214e-10, 2.062158e-10, 
    2.071446e-10, 2.073314e-10, 2.059205e-10, 2.067861e-10, 2.040154e-10, 
    2.044616e-10, 2.041959e-10, 2.032269e-10, 2.063322e-10, 2.047352e-10, 
    2.076898e-10, 2.068205e-10, 2.093635e-10, 2.080966e-10, 2.105892e-10, 
    2.1166e-10, 2.126708e-10, 2.138555e-10, 2.039541e-10, 2.036171e-10, 
    2.042208e-10, 2.050577e-10, 2.058361e-10, 2.068734e-10, 2.069798e-10, 
    2.071745e-10, 2.076794e-10, 2.081045e-10, 2.072361e-10, 2.082111e-10, 
    2.045651e-10, 2.064712e-10, 2.034897e-10, 2.043849e-10, 2.050084e-10, 
    2.047347e-10, 2.06158e-10, 2.064943e-10, 2.078641e-10, 2.071554e-10, 
    2.113954e-10, 2.095134e-10, 2.147602e-10, 2.132863e-10, 2.034994e-10, 
    2.03953e-10, 2.05536e-10, 2.04782e-10, 2.069428e-10, 2.074767e-10, 
    2.079113e-10, 2.084676e-10, 2.085278e-10, 2.088578e-10, 2.083171e-10, 
    2.088364e-10, 2.068757e-10, 2.077506e-10, 2.053548e-10, 2.059364e-10, 
    2.056687e-10, 2.053753e-10, 2.062817e-10, 2.072497e-10, 2.072705e-10, 
    2.075815e-10, 2.084592e-10, 2.069516e-10, 2.11639e-10, 2.08737e-10, 
    2.044482e-10, 2.053247e-10, 2.054501e-10, 2.051102e-10, 2.074231e-10, 
    2.065834e-10, 2.088498e-10, 2.082358e-10, 2.092423e-10, 2.087418e-10, 
    2.086682e-10, 2.080266e-10, 2.076277e-10, 2.066218e-10, 2.058055e-10, 
    2.051595e-10, 2.053096e-10, 2.060196e-10, 2.073091e-10, 2.085332e-10, 
    2.082647e-10, 2.091657e-10, 2.067857e-10, 2.077818e-10, 2.073965e-10, 
    2.08402e-10, 2.062024e-10, 2.080745e-10, 2.057254e-10, 2.059307e-10, 
    2.065667e-10, 2.078494e-10, 2.081339e-10, 2.084378e-10, 2.082502e-10, 
    2.073419e-10, 2.071932e-10, 2.065512e-10, 2.063742e-10, 2.05886e-10, 
    2.054823e-10, 2.058511e-10, 2.062388e-10, 2.073422e-10, 2.083395e-10, 
    2.094299e-10, 2.096973e-10, 2.109764e-10, 2.099348e-10, 2.116552e-10, 
    2.10192e-10, 2.127288e-10, 2.081834e-10, 2.10149e-10, 2.065957e-10, 
    2.069768e-10, 2.076672e-10, 2.092557e-10, 2.083973e-10, 2.094014e-10, 
    2.071874e-10, 2.060441e-10, 2.057489e-10, 2.051987e-10, 2.057614e-10, 
    2.057157e-10, 2.062549e-10, 2.060815e-10, 2.073789e-10, 2.066814e-10, 
    2.086664e-10, 2.093935e-10, 2.114547e-10, 2.127241e-10, 2.140209e-10, 
    2.145949e-10, 2.147697e-10, 2.148429e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24786.37, 24802.16, 24799.07, 24811.95, 24804.78, 24813.24, 24789.55, 
    24802.79, 24794.32, 24787.78, 24837.42, 24812.53, 24863.9, 24847.59, 
    24889.18, 24861.34, 24894.84, 24888.36, 24907.92, 24902.28, 24927.75, 
    24910.53, 24941.27, 24923.61, 24926.35, 24909.97, 24817.48, 24834.28, 
    24816.49, 24818.87, 24817.8, 24804.93, 24798.5, 24785.17, 24787.58, 
    24797.38, 24819.94, 24812.23, 24831.78, 24831.34, 24853.56, 24843.5, 
    24881.56, 24870.57, 24902.51, 24894.45, 24902.13, 24899.79, 24902.16, 
    24890.36, 24895.4, 24885, 24845.38, 24856.85, 24822.95, 24803.1, 
    24790.13, 24781.02, 24782.3, 24784.75, 24797.43, 24809.51, 24818.79, 
    24825.06, 24831.27, 24850.33, 24860.52, 24883.79, 24879.55, 24886.76, 
    24893.65, 24905.25, 24903.33, 24908.48, 24886.56, 24901.09, 24877.14, 
    24883.67, 24832.98, 24814.3, 24806.47, 24799.66, 24783.29, 24794.57, 
    24790.11, 24800.75, 24807.58, 24804.19, 24825.23, 24817, 24861.13, 
    24841.91, 24892.85, 24880.42, 24895.82, 24887.96, 24901.44, 24889.32, 
    24910.4, 24915.06, 24911.87, 24924.17, 24888.64, 24902.13, 24804.1, 
    24804.65, 24807.22, 24795.98, 24795.29, 24785.11, 24794.17, 24798.05, 
    24807.97, 24813.89, 24819.54, 24832.09, 24846.31, 24866.46, 24881.22, 
    24891.26, 24885.09, 24890.54, 24884.45, 24881.61, 24913.31, 24895.45, 
    24922.39, 24920.88, 24908.6, 24921.05, 24805.04, 24801.87, 24790.96, 
    24799.49, 24784, 24792.64, 24797.64, 24817.17, 24821.51, 24825.55, 
    24833.59, 24844.01, 24862.49, 24878.87, 24894.05, 24892.95, 24893.33, 
    24896.72, 24888.32, 24898.1, 24899.74, 24895.45, 24920.67, 24913.39, 
    24920.85, 24916.09, 24802.9, 24808.24, 24805.35, 24810.79, 24806.95, 
    24824.1, 24829.3, 24854, 24843.81, 24860.07, 24845.45, 24848.04, 
    24860.61, 24846.24, 24877.96, 24856.34, 24896.85, 24874.88, 24898.23, 
    24893.99, 24901.02, 24907.37, 24915.43, 24930.51, 24926.99, 24939.77, 
    24816.24, 24823.26, 24822.63, 24830.03, 24835.54, 24847.59, 24867.14, 
    24859.73, 24873.37, 24876.14, 24855.43, 24868.09, 24827.98, 24834.37, 
    24830.56, 24816.79, 24861.44, 24838.3, 24881.47, 24868.59, 24906.46, 
    24887.55, 24925.06, 24941.62, 24957.5, 24976.49, 24827.11, 24822.31, 
    24830.91, 24842.95, 24854.21, 24869.37, 24870.94, 24873.82, 24881.31, 
    24887.66, 24874.73, 24889.26, 24835.86, 24863.47, 24820.51, 24833.27, 
    24842.24, 24838.29, 24858.89, 24863.8, 24884.07, 24873.53, 24937.5, 
    24908.72, 24991.25, 24967.32, 24820.64, 24827.09, 24849.87, 24838.97, 
    24870.39, 24878.29, 24884.77, 24893.09, 24893.98, 24898.89, 24890.86, 
    24898.57, 24869.41, 24882.37, 24847.25, 24855.67, 24851.78, 24847.54, 
    24860.7, 24874.93, 24875.24, 24879.85, 24892.97, 24870.52, 24941.29, 
    24897.1, 24834.17, 24846.81, 24848.62, 24843.71, 24877.5, 24865.11, 
    24898.77, 24889.63, 24904.64, 24897.16, 24896.07, 24886.5, 24880.54, 
    24865.68, 24853.77, 24844.42, 24846.59, 24856.88, 24875.81, 24894.06, 
    24890.07, 24903.49, 24868.08, 24882.84, 24877.11, 24892.12, 24859.54, 
    24887.22, 24852.6, 24855.58, 24864.87, 24883.85, 24888.1, 24892.65, 
    24889.85, 24876.29, 24874.09, 24864.64, 24862.05, 24854.93, 24849.09, 
    24854.43, 24860.07, 24876.3, 24891.19, 24907.46, 24911.49, 24931.02, 
    24915.09, 24941.55, 24919.01, 24958.43, 24888.85, 24918.35, 24865.29, 
    24870.9, 24881.13, 24904.85, 24892.04, 24907.04, 24874.01, 24857.23, 
    24852.95, 24844.99, 24853.13, 24852.46, 24860.3, 24857.78, 24876.84, 
    24866.55, 24896.04, 24906.92, 24938.42, 24958.35, 24979.16, 24988.53, 
    24991.4, 24992.61 ;

 GC_ICE1 =
  17951.62, 17976.51, 17971.64, 17991.95, 17980.65, 17993.99, 17956.64, 
    17977.51, 17964.16, 17953.85, 18032.07, 17992.86, 18073.76, 18048.08, 
    18113.52, 18069.73, 18122.41, 18112.23, 18142.93, 18134.09, 18174.06, 
    18147.03, 18195.27, 18167.55, 18171.85, 18146.15, 18000.66, 18027.13, 
    17999.11, 18002.85, 18001.17, 17980.88, 17970.75, 17949.74, 17953.53, 
    17968.98, 18004.53, 17992.39, 18023.2, 18022.49, 18057.49, 18041.65, 
    18101.53, 18084.25, 18134.45, 18121.8, 18133.86, 18130.19, 18133.9, 
    18115.38, 18123.3, 18106.95, 18044.62, 18062.66, 18009.28, 17978.01, 
    17957.55, 17943.19, 17945.21, 17949.08, 17969.07, 17988.1, 18002.73, 
    18012.6, 18022.39, 18052.4, 18068.44, 18105.05, 18098.37, 18109.71, 
    18120.55, 18138.74, 18135.73, 18143.81, 18109.41, 18132.22, 18094.58, 
    18104.85, 18025.07, 17995.65, 17983.32, 17972.58, 17946.77, 17964.55, 
    17957.52, 17974.29, 17985.05, 17979.72, 18012.87, 17999.91, 18069.4, 
    18039.15, 18119.3, 18099.74, 18123.95, 18111.61, 18132.76, 18113.74, 
    18146.83, 18154.14, 18149.14, 18168.44, 18112.68, 18133.86, 17979.57, 
    17980.44, 17984.49, 17966.77, 17965.7, 17949.63, 17963.92, 17970.04, 
    17985.68, 17995, 18003.9, 18023.67, 18046.07, 18077.78, 18101, 18116.79, 
    18107.09, 18115.66, 18106.08, 18101.62, 18151.39, 18123.37, 18165.64, 
    18163.27, 18144, 18163.54, 17981.05, 17976.06, 17958.86, 17972.31, 
    17947.89, 17961.52, 17969.4, 18000.18, 18007.01, 18013.38, 18026.04, 
    18042.46, 18071.53, 18097.3, 18121.18, 18119.44, 18120.05, 18125.36, 
    18112.17, 18127.52, 18130.11, 18123.37, 18162.95, 18151.52, 18163.22, 
    18155.76, 17977.68, 17986.1, 17981.54, 17990.12, 17984.07, 18011.09, 
    18019.29, 18058.17, 18042.14, 18067.72, 18044.73, 18048.79, 18068.57, 
    18045.97, 18095.87, 18061.85, 18125.57, 18091.02, 18127.73, 18121.07, 
    18132.11, 18142.08, 18154.72, 18178.38, 18172.87, 18192.9, 17998.71, 
    18009.76, 18008.78, 18020.43, 18029.11, 18048.09, 18078.85, 18067.2, 
    18088.66, 18093.01, 18060.43, 18080.34, 18017.21, 18027.26, 18021.26, 
    17999.58, 18069.88, 18033.46, 18101.39, 18081.14, 18140.65, 18110.96, 
    18169.84, 18195.81, 18220.73, 18250.5, 18015.83, 18008.28, 18021.82, 
    18040.79, 18058.51, 18082.37, 18084.83, 18089.35, 18101.14, 18111.14, 
    18090.79, 18113.65, 18029.61, 18073.07, 18005.43, 18025.53, 18039.66, 
    18033.44, 18065.87, 18073.61, 18105.48, 18088.91, 18189.35, 18144.2, 
    18273.64, 18236.12, 18005.65, 18015.8, 18051.67, 18034.52, 18083.97, 
    18096.4, 18106.59, 18119.67, 18121.06, 18128.77, 18116.16, 18128.27, 
    18082.42, 18102.81, 18047.55, 18060.8, 18054.69, 18048.02, 18068.71, 
    18091.11, 18091.59, 18098.85, 18119.48, 18084.18, 18195.3, 18125.96, 
    18026.96, 18046.87, 18049.72, 18041.98, 18095.15, 18075.66, 18128.58, 
    18114.24, 18137.79, 18126.06, 18124.34, 18109.3, 18099.93, 18076.55, 
    18057.81, 18043.1, 18046.52, 18062.7, 18092.49, 18121.19, 18114.92, 
    18135.99, 18080.33, 18103.55, 18094.53, 18118.14, 18066.89, 18110.45, 
    18055.98, 18060.67, 18075.27, 18105.14, 18111.83, 18118.97, 18114.58, 
    18093.25, 18089.79, 18074.92, 18070.84, 18059.65, 18050.45, 18058.85, 
    18067.73, 18093.26, 18116.69, 18142.22, 18148.54, 18179.18, 18154.19, 
    18195.7, 18160.33, 18222.18, 18113.01, 18159.3, 18075.94, 18084.76, 
    18100.86, 18138.12, 18118.03, 18141.55, 18089.65, 18063.27, 18056.52, 
    18043.99, 18056.8, 18055.76, 18068.1, 18064.12, 18094.12, 18077.92, 
    18124.3, 18141.36, 18190.79, 18222.06, 18254.7, 18269.38, 18273.89, 
    18275.78 ;

 GC_LIQ1 =
  5291.727, 5293.509, 5293.16, 5294.615, 5293.805, 5294.762, 5292.086, 
    5293.58, 5292.624, 5291.886, 5297.501, 5294.68, 5300.52, 5298.655, 
    5303.409, 5300.228, 5304.064, 5303.316, 5305.585, 5304.93, 5307.894, 
    5305.89, 5309.469, 5307.411, 5307.73, 5305.824, 5295.242, 5297.146, 
    5295.13, 5295.399, 5295.278, 5293.822, 5293.096, 5291.592, 5291.864, 
    5292.969, 5295.52, 5294.646, 5296.863, 5296.812, 5299.338, 5298.191, 
    5302.538, 5301.282, 5304.957, 5304.019, 5304.913, 5304.641, 5304.916, 
    5303.545, 5304.13, 5302.932, 5298.405, 5299.713, 5295.861, 5293.616, 
    5292.151, 5291.125, 5291.269, 5291.545, 5292.975, 5294.339, 5295.391, 
    5296.1, 5296.805, 5298.969, 5300.133, 5302.794, 5302.308, 5303.132, 
    5303.926, 5305.275, 5305.052, 5305.65, 5303.11, 5304.791, 5302.033, 
    5302.779, 5296.998, 5294.881, 5293.996, 5293.227, 5291.38, 5292.652, 
    5292.148, 5293.35, 5294.121, 5293.739, 5296.12, 5295.188, 5300.203, 
    5298.011, 5303.833, 5302.408, 5304.179, 5303.271, 5304.832, 5303.426, 
    5305.875, 5306.417, 5306.045, 5307.477, 5303.348, 5304.913, 5293.728, 
    5293.79, 5294.081, 5292.811, 5292.734, 5291.585, 5292.606, 5293.044, 
    5294.166, 5294.834, 5295.475, 5296.897, 5298.51, 5300.812, 5302.5, 
    5303.648, 5302.942, 5303.565, 5302.869, 5302.544, 5306.213, 5304.135, 
    5307.27, 5307.094, 5305.665, 5307.114, 5293.834, 5293.476, 5292.245, 
    5293.208, 5291.46, 5292.435, 5292.999, 5295.207, 5295.698, 5296.157, 
    5297.067, 5298.25, 5300.358, 5302.23, 5303.973, 5303.844, 5303.89, 
    5304.283, 5303.312, 5304.443, 5304.634, 5304.135, 5307.07, 5306.222, 
    5307.09, 5306.537, 5293.592, 5294.195, 5293.869, 5294.483, 5294.05, 
    5295.992, 5296.581, 5299.388, 5298.226, 5300.082, 5298.413, 5298.707, 
    5300.143, 5298.502, 5302.126, 5299.655, 5304.298, 5301.774, 5304.458, 
    5303.965, 5304.783, 5305.522, 5306.459, 5308.215, 5307.806, 5309.293, 
    5295.101, 5295.896, 5295.826, 5296.664, 5297.289, 5298.656, 5300.89, 
    5300.043, 5301.603, 5301.918, 5299.552, 5300.998, 5296.432, 5297.155, 
    5296.724, 5295.164, 5300.238, 5297.601, 5302.528, 5301.056, 5305.417, 
    5303.223, 5307.581, 5309.509, 5311.36, 5313.573, 5296.333, 5295.79, 
    5296.764, 5298.129, 5299.412, 5301.145, 5301.324, 5301.653, 5302.51, 
    5303.236, 5301.757, 5303.419, 5297.324, 5300.47, 5295.585, 5297.031, 
    5298.048, 5297.6, 5299.947, 5300.509, 5302.825, 5301.621, 5309.029, 
    5305.679, 5315.295, 5312.504, 5295.6, 5296.331, 5298.916, 5297.677, 
    5301.262, 5302.165, 5302.906, 5303.861, 5303.964, 5304.536, 5303.602, 
    5304.499, 5301.149, 5302.631, 5298.617, 5299.579, 5299.135, 5298.65, 
    5300.153, 5301.78, 5301.815, 5302.343, 5303.847, 5301.277, 5309.471, 
    5304.327, 5297.133, 5298.567, 5298.774, 5298.214, 5302.074, 5300.658, 
    5304.521, 5303.462, 5305.205, 5304.334, 5304.207, 5303.103, 5302.422, 
    5300.722, 5299.361, 5298.295, 5298.542, 5299.717, 5301.881, 5303.974, 
    5303.512, 5305.071, 5300.998, 5302.685, 5302.029, 5303.748, 5300.021, 
    5303.186, 5299.229, 5299.569, 5300.63, 5302.8, 5303.287, 5303.81, 
    5303.486, 5301.937, 5301.685, 5300.604, 5300.308, 5299.495, 5298.827, 
    5299.437, 5300.082, 5301.937, 5303.64, 5305.533, 5306.001, 5308.274, 
    5306.42, 5309.5, 5306.876, 5311.468, 5303.372, 5306.799, 5300.678, 
    5301.319, 5302.489, 5305.229, 5303.74, 5305.483, 5301.675, 5299.758, 
    5299.268, 5298.36, 5299.289, 5299.212, 5300.108, 5299.82, 5301.999, 
    5300.822, 5304.204, 5305.469, 5309.136, 5311.459, 5313.885, 5314.978, 
    5315.313, 5315.454 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  1.074026e-08, 1.076965e-08, 1.076394e-08, 1.078764e-08, 1.07745e-08, 
    1.079002e-08, 1.074622e-08, 1.077082e-08, 1.075512e-08, 1.074291e-08, 
    1.083362e-08, 1.07887e-08, 1.088028e-08, 1.085164e-08, 1.092357e-08, 
    1.087582e-08, 1.09332e-08, 1.09222e-08, 1.095531e-08, 1.094583e-08, 
    1.098816e-08, 1.095969e-08, 1.10101e-08, 1.098136e-08, 1.098586e-08, 
    1.095875e-08, 1.079775e-08, 1.082803e-08, 1.079595e-08, 1.080027e-08, 
    1.079833e-08, 1.077477e-08, 1.076289e-08, 1.073801e-08, 1.074253e-08, 
    1.07608e-08, 1.080221e-08, 1.078816e-08, 1.082358e-08, 1.082278e-08, 
    1.08622e-08, 1.084443e-08, 1.091066e-08, 1.089184e-08, 1.094622e-08, 
    1.093255e-08, 1.094558e-08, 1.094163e-08, 1.094563e-08, 1.092558e-08, 
    1.093417e-08, 1.091652e-08, 1.084776e-08, 1.086797e-08, 1.080767e-08, 
    1.077139e-08, 1.07473e-08, 1.07302e-08, 1.073261e-08, 1.073722e-08, 
    1.076091e-08, 1.078318e-08, 1.080014e-08, 1.081149e-08, 1.082267e-08, 
    1.085649e-08, 1.087439e-08, 1.091447e-08, 1.090724e-08, 1.091949e-08, 
    1.093119e-08, 1.095083e-08, 1.09476e-08, 1.095625e-08, 1.091917e-08, 
    1.094381e-08, 1.090312e-08, 1.091425e-08, 1.082569e-08, 1.079195e-08, 
    1.077759e-08, 1.076504e-08, 1.073447e-08, 1.075558e-08, 1.074726e-08, 
    1.076706e-08, 1.077963e-08, 1.077342e-08, 1.08118e-08, 1.079688e-08, 
    1.087545e-08, 1.084161e-08, 1.092982e-08, 1.090872e-08, 1.093488e-08, 
    1.092154e-08, 1.09444e-08, 1.092382e-08, 1.095947e-08, 1.096723e-08, 
    1.096193e-08, 1.09823e-08, 1.092268e-08, 1.094558e-08, 1.077324e-08, 
    1.077425e-08, 1.077898e-08, 1.07582e-08, 1.075693e-08, 1.073789e-08, 
    1.075483e-08, 1.076205e-08, 1.078036e-08, 1.079119e-08, 1.080149e-08, 
    1.082412e-08, 1.084939e-08, 1.088472e-08, 1.091009e-08, 1.09271e-08, 
    1.091667e-08, 1.092588e-08, 1.091558e-08, 1.091076e-08, 1.096432e-08, 
    1.093425e-08, 1.097937e-08, 1.097687e-08, 1.095645e-08, 1.097716e-08, 
    1.077497e-08, 1.076913e-08, 1.074886e-08, 1.076472e-08, 1.073582e-08, 
    1.0752e-08, 1.07613e-08, 1.079718e-08, 1.080507e-08, 1.081238e-08, 
    1.082682e-08, 1.084534e-08, 1.087782e-08, 1.090608e-08, 1.093187e-08, 
    1.092998e-08, 1.093065e-08, 1.093641e-08, 1.092214e-08, 1.093875e-08, 
    1.094153e-08, 1.093425e-08, 1.097654e-08, 1.096446e-08, 1.097682e-08, 
    1.096896e-08, 1.077103e-08, 1.078085e-08, 1.077554e-08, 1.078552e-08, 
    1.077849e-08, 1.080975e-08, 1.081912e-08, 1.086296e-08, 1.084497e-08, 
    1.08736e-08, 1.084788e-08, 1.085244e-08, 1.087453e-08, 1.084927e-08, 
    1.090452e-08, 1.086706e-08, 1.093663e-08, 1.089923e-08, 1.093897e-08, 
    1.093176e-08, 1.09437e-08, 1.09544e-08, 1.096785e-08, 1.099267e-08, 
    1.098693e-08, 1.100768e-08, 1.079549e-08, 1.080823e-08, 1.080711e-08, 
    1.082044e-08, 1.083029e-08, 1.085165e-08, 1.08859e-08, 1.087302e-08, 
    1.089666e-08, 1.090141e-08, 1.086549e-08, 1.088754e-08, 1.081675e-08, 
    1.082819e-08, 1.082138e-08, 1.079649e-08, 1.087599e-08, 1.08352e-08, 
    1.091051e-08, 1.088842e-08, 1.095287e-08, 1.092082e-08, 1.098376e-08, 
    1.101065e-08, 1.103597e-08, 1.106552e-08, 1.081518e-08, 1.080653e-08, 
    1.082202e-08, 1.084345e-08, 1.086334e-08, 1.088977e-08, 1.089247e-08, 
    1.089742e-08, 1.091025e-08, 1.092103e-08, 1.089899e-08, 1.092373e-08, 
    1.083084e-08, 1.087953e-08, 1.080325e-08, 1.082622e-08, 1.084219e-08, 
    1.083519e-08, 1.087155e-08, 1.088012e-08, 1.091493e-08, 1.089694e-08, 
    1.100401e-08, 1.095665e-08, 1.108803e-08, 1.105133e-08, 1.08035e-08, 
    1.081515e-08, 1.085568e-08, 1.08364e-08, 1.089153e-08, 1.09051e-08, 
    1.091613e-08, 1.093022e-08, 1.093175e-08, 1.09401e-08, 1.092641e-08, 
    1.093956e-08, 1.088983e-08, 1.091205e-08, 1.085105e-08, 1.08659e-08, 
    1.085907e-08, 1.085157e-08, 1.08747e-08, 1.089933e-08, 1.089986e-08, 
    1.090776e-08, 1.093e-08, 1.089176e-08, 1.101011e-08, 1.093703e-08, 
    1.082785e-08, 1.085028e-08, 1.085348e-08, 1.08448e-08, 1.090374e-08, 
    1.088239e-08, 1.093989e-08, 1.092435e-08, 1.094981e-08, 1.093716e-08, 
    1.09353e-08, 1.091905e-08, 1.090893e-08, 1.088336e-08, 1.086256e-08, 
    1.084606e-08, 1.084989e-08, 1.086802e-08, 1.090084e-08, 1.093188e-08, 
    1.092508e-08, 1.094788e-08, 1.088754e-08, 1.091284e-08, 1.090306e-08, 
    1.092856e-08, 1.087268e-08, 1.092025e-08, 1.086051e-08, 1.086576e-08, 
    1.088196e-08, 1.091455e-08, 1.092177e-08, 1.092947e-08, 1.092472e-08, 
    1.090167e-08, 1.08979e-08, 1.088157e-08, 1.087706e-08, 1.086461e-08, 
    1.085431e-08, 1.086372e-08, 1.087361e-08, 1.090168e-08, 1.092698e-08, 
    1.095455e-08, 1.09613e-08, 1.099349e-08, 1.096728e-08, 1.101052e-08, 
    1.097375e-08, 1.10374e-08, 1.092302e-08, 1.097267e-08, 1.08827e-08, 
    1.08924e-08, 1.090993e-08, 1.095015e-08, 1.092844e-08, 1.095383e-08, 
    1.089775e-08, 1.086864e-08, 1.086111e-08, 1.084706e-08, 1.086144e-08, 
    1.086027e-08, 1.087402e-08, 1.08696e-08, 1.090262e-08, 1.088488e-08, 
    1.093525e-08, 1.095363e-08, 1.100551e-08, 1.103729e-08, 1.106965e-08, 
    1.108393e-08, 1.108827e-08, 1.109009e-08 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.431473, 6.459629, 6.454149, 6.476902, 6.464273, 6.479182, 6.437174, 
    6.46075, 6.445693, 6.434003, 6.521199, 6.477918, 6.566323, 6.538589, 
    6.608384, 6.562005, 6.617757, 6.607039, 6.63932, 6.630063, 6.671458, 
    6.643595, 6.692968, 6.664796, 6.6692, 6.642677, 6.486611, 6.515802, 
    6.484885, 6.489042, 6.487175, 6.464535, 6.453146, 6.429322, 6.433643, 
    6.451141, 6.490911, 6.477393, 6.511489, 6.510717, 6.548801, 6.531614, 
    6.595817, 6.577531, 6.630449, 6.617118, 6.629823, 6.625968, 6.629873, 
    6.610328, 6.618698, 6.601513, 6.534832, 6.554389, 6.496163, 6.461306, 
    6.438208, 6.421849, 6.42416, 6.428568, 6.451244, 6.472604, 6.488912, 
    6.499835, 6.510607, 6.543287, 6.560616, 6.59952, 6.592486, 6.604402, 
    6.615793, 6.634946, 6.631791, 6.640238, 6.604085, 6.628101, 6.588482, 
    6.599305, 6.513549, 6.481038, 6.467258, 6.455203, 6.425938, 6.446139, 
    6.438171, 6.457135, 6.469203, 6.463233, 6.500133, 6.485773, 6.561644, 
    6.5289, 6.614463, 6.593929, 6.61939, 6.60639, 6.628675, 6.608617, 
    6.643383, 6.650969, 6.645784, 6.665707, 6.607506, 6.629824, 6.463066, 
    6.464039, 6.468575, 6.448651, 6.447433, 6.429204, 6.445421, 6.452335, 
    6.469903, 6.480309, 6.490211, 6.512012, 6.536413, 6.570621, 6.595259, 
    6.611805, 6.601655, 6.610616, 6.6006, 6.595909, 6.648127, 6.618777, 
    6.662839, 6.660396, 6.64044, 6.660671, 6.464723, 6.459121, 6.439698, 
    6.454895, 6.427221, 6.442704, 6.451618, 6.486075, 6.493658, 6.500697, 
    6.51461, 6.532493, 6.563935, 6.591362, 6.616455, 6.614614, 6.615263, 
    6.620876, 6.606977, 6.62316, 6.625879, 6.618772, 6.660069, 6.648256, 
    6.660344, 6.65265, 6.460941, 6.47037, 6.465274, 6.474859, 6.468107, 
    6.498168, 6.507197, 6.549542, 6.532141, 6.559845, 6.534951, 6.539359, 
    6.560755, 6.536294, 6.58985, 6.553517, 6.621095, 6.584718, 6.623378, 
    6.616346, 6.62799, 6.63843, 6.651575, 6.675871, 6.67024, 6.690586, 
    6.484441, 6.496699, 6.495617, 6.508458, 6.517965, 6.538595, 6.571767, 
    6.55928, 6.582211, 6.586821, 6.551987, 6.573364, 6.50491, 6.515943, 
    6.509371, 6.485408, 6.56216, 6.522705, 6.595667, 6.574212, 6.636941, 
    6.605704, 6.667142, 6.693511, 6.718372, 6.747504, 6.503393, 6.495057, 
    6.509985, 6.530677, 6.549904, 6.57552, 6.578143, 6.58295, 6.595408, 
    6.605896, 6.584473, 6.608525, 6.518508, 6.56559, 6.49191, 6.514048, 
    6.529455, 6.522691, 6.557854, 6.566158, 6.599968, 6.582476, 6.687, 
    6.640639, 6.769724, 6.733511, 6.492146, 6.503363, 6.542494, 6.523858, 
    6.577231, 6.590408, 6.60113, 6.614854, 6.616335, 6.624475, 6.61114, 
    6.623948, 6.575574, 6.597166, 6.538011, 6.552382, 6.545768, 6.538519, 
    6.560906, 6.58481, 6.585318, 6.592994, 6.614661, 6.577447, 6.693004, 
    6.621509, 6.515608, 6.537274, 6.540368, 6.531968, 6.589087, 6.568357, 
    6.624276, 6.609136, 6.633953, 6.621614, 6.619801, 6.603974, 6.594133, 
    6.569308, 6.549148, 6.533185, 6.536895, 6.554436, 6.586273, 6.616471, 
    6.60985, 6.632065, 6.573352, 6.597937, 6.588429, 6.613235, 6.558949, 
    6.605172, 6.547167, 6.55224, 6.567946, 6.599609, 6.60662, 6.614118, 
    6.60949, 6.587082, 6.583413, 6.567564, 6.563193, 6.551135, 6.541163, 
    6.550274, 6.559852, 6.58709, 6.611694, 6.638579, 6.645166, 6.676685, 
    6.651026, 6.693404, 6.657373, 6.71981, 6.60785, 6.656308, 6.56866, 
    6.57807, 6.595112, 6.634289, 6.613118, 6.637879, 6.583269, 6.555044, 
    6.547748, 6.534156, 6.548059, 6.546927, 6.560246, 6.555964, 6.587995, 
    6.570778, 6.619756, 6.637682, 6.688453, 6.719688, 6.751562, 6.765662, 
    6.769957, 6.771753,
  4.809054, 4.826082, 4.822768, 4.836523, 4.828888, 4.837901, 4.812501, 
    4.82676, 4.817654, 4.810583, 4.863285, 4.837137, 4.890507, 4.873774, 
    4.915859, 4.887904, 4.921505, 4.915046, 4.934487, 4.928913, 4.953834, 
    4.937061, 4.96677, 4.949823, 4.952474, 4.936509, 4.842388, 4.860027, 
    4.841345, 4.843858, 4.842729, 4.829048, 4.822164, 4.807751, 4.810365, 
    4.82095, 4.844988, 4.836817, 4.857413, 4.856947, 4.879935, 4.869563, 
    4.908284, 4.897261, 4.929146, 4.921118, 4.92877, 4.926448, 4.9288, 
    4.917028, 4.92207, 4.911716, 4.871506, 4.883307, 4.848159, 4.8271, 
    4.813128, 4.80323, 4.804628, 4.807296, 4.821012, 4.833923, 4.843777, 
    4.850375, 4.856881, 4.876614, 4.887064, 4.910517, 4.906276, 4.913458, 
    4.920319, 4.931855, 4.929955, 4.935041, 4.913266, 4.927734, 4.903862, 
    4.910386, 4.858667, 4.83902, 4.830697, 4.823405, 4.805704, 4.817925, 
    4.813106, 4.824572, 4.831868, 4.828259, 4.850556, 4.841881, 4.887684, 
    4.867927, 4.919518, 4.907146, 4.922486, 4.914654, 4.928079, 4.915996, 
    4.936934, 4.941501, 4.93838, 4.950369, 4.915327, 4.928771, 4.828158, 
    4.828747, 4.831488, 4.819444, 4.818707, 4.80768, 4.81749, 4.821671, 
    4.83229, 4.83858, 4.844563, 4.85773, 4.872461, 4.893096, 4.907948, 
    4.917917, 4.911801, 4.9172, 4.911166, 4.908338, 4.939791, 4.922118, 
    4.948644, 4.947174, 4.935163, 4.947339, 4.82916, 4.825773, 4.814028, 
    4.823218, 4.80648, 4.815847, 4.821239, 4.842066, 4.846644, 4.850897, 
    4.859298, 4.870094, 4.889064, 4.9056, 4.920718, 4.919609, 4.919999, 
    4.923381, 4.915009, 4.924757, 4.926395, 4.922114, 4.946977, 4.939867, 
    4.947142, 4.942512, 4.826873, 4.832573, 4.829493, 4.835287, 4.831206, 
    4.849372, 4.854826, 4.880385, 4.869882, 4.886598, 4.871578, 4.874238, 
    4.887151, 4.872387, 4.90469, 4.882784, 4.923513, 4.901599, 4.924888, 
    4.920652, 4.927665, 4.933952, 4.941864, 4.956486, 4.953098, 4.965335, 
    4.841076, 4.848484, 4.847828, 4.855584, 4.861324, 4.873776, 4.893786, 
    4.886255, 4.900082, 4.902862, 4.881855, 4.89475, 4.853442, 4.860106, 
    4.856135, 4.841662, 4.887995, 4.864189, 4.908194, 4.89526, 4.933056, 
    4.914244, 4.951233, 4.967099, 4.982039, 4.999546, 4.852525, 4.847489, 
    4.856505, 4.869, 4.8806, 4.896049, 4.89763, 4.900528, 4.908037, 4.914356, 
    4.901448, 4.915941, 4.861659, 4.890063, 4.845589, 4.858963, 4.868262, 
    4.864178, 4.885394, 4.890403, 4.910787, 4.900242, 4.963184, 4.935285, 
    5.012886, 4.991139, 4.845731, 4.852507, 4.876131, 4.864882, 4.89708, 
    4.905024, 4.911485, 4.919755, 4.920646, 4.92555, 4.917516, 4.925231, 
    4.896082, 4.909096, 4.873423, 4.882095, 4.878103, 4.87373, 4.887236, 
    4.901652, 4.901955, 4.906584, 4.919648, 4.897211, 4.9668, 4.923772, 
    4.8599, 4.872983, 4.874846, 4.869776, 4.904228, 4.89173, 4.925429, 
    4.916308, 4.931256, 4.923826, 4.922733, 4.913199, 4.907269, 4.892304, 
    4.880144, 4.870511, 4.87275, 4.883335, 4.902534, 4.920729, 4.916741, 
    4.930119, 4.894742, 4.909563, 4.903833, 4.918778, 4.886056, 4.913929, 
    4.878947, 4.882008, 4.891482, 4.910572, 4.914793, 4.919312, 4.916522, 
    4.90302, 4.900808, 4.891251, 4.888617, 4.881341, 4.875325, 4.880823, 
    4.886601, 4.903024, 4.917851, 4.934042, 4.938007, 4.956981, 4.94154, 
    4.967041, 4.945367, 4.982912, 4.91554, 4.944719, 4.891912, 4.897585, 
    4.907862, 4.931462, 4.918708, 4.933623, 4.900721, 4.883703, 4.879298, 
    4.871097, 4.879486, 4.878803, 4.886837, 4.884254, 4.90357, 4.893189, 
    4.922707, 4.933504, 4.964054, 4.982834, 5.001979, 5.010446, 5.013024, 
    5.014102,
  4.269382, 4.283989, 4.281146, 4.292946, 4.286397, 4.294128, 4.272339, 
    4.284571, 4.276759, 4.270693, 4.315906, 4.293473, 4.339261, 4.324905, 
    4.361014, 4.337028, 4.365859, 4.360317, 4.376999, 4.372216, 4.393601, 
    4.379208, 4.404703, 4.390159, 4.392434, 4.378734, 4.297978, 4.31311, 
    4.297083, 4.299239, 4.298271, 4.286533, 4.280628, 4.268264, 4.270506, 
    4.279587, 4.300208, 4.293199, 4.310869, 4.310469, 4.330191, 4.321292, 
    4.354515, 4.345057, 4.372416, 4.365527, 4.372093, 4.3701, 4.372118, 
    4.362017, 4.366344, 4.35746, 4.322959, 4.333084, 4.302929, 4.284862, 
    4.272876, 4.264386, 4.265585, 4.267874, 4.27964, 4.290717, 4.29917, 
    4.304831, 4.310411, 4.327341, 4.336308, 4.356431, 4.352792, 4.358954, 
    4.364841, 4.37474, 4.37311, 4.377475, 4.358789, 4.371204, 4.35072, 
    4.356318, 4.311944, 4.295089, 4.287948, 4.281693, 4.266508, 4.276992, 
    4.272858, 4.282694, 4.288953, 4.285857, 4.304986, 4.297543, 4.33684, 
    4.319888, 4.364155, 4.353538, 4.366701, 4.359981, 4.3715, 4.361132, 
    4.379098, 4.383018, 4.38034, 4.390628, 4.360558, 4.372094, 4.28577, 
    4.286275, 4.288627, 4.278295, 4.277663, 4.268203, 4.276618, 4.280206, 
    4.289315, 4.294712, 4.299844, 4.31114, 4.323779, 4.341483, 4.354226, 
    4.36278, 4.357533, 4.362165, 4.356987, 4.354561, 4.38155, 4.366385, 
    4.389147, 4.387886, 4.377579, 4.388028, 4.28663, 4.283724, 4.273649, 
    4.281533, 4.267174, 4.275209, 4.279835, 4.297702, 4.30163, 4.305278, 
    4.312486, 4.321748, 4.338024, 4.352211, 4.365183, 4.364232, 4.364567, 
    4.367469, 4.360284, 4.368649, 4.370055, 4.366382, 4.387717, 4.381615, 
    4.387859, 4.383885, 4.284668, 4.289558, 4.286916, 4.291886, 4.288385, 
    4.303969, 4.308648, 4.330577, 4.321566, 4.335907, 4.32302, 4.325304, 
    4.336382, 4.323716, 4.351431, 4.332635, 4.367582, 4.348778, 4.368762, 
    4.365128, 4.371145, 4.37654, 4.38333, 4.395877, 4.39297, 4.403472, 
    4.296853, 4.303207, 4.302645, 4.309299, 4.314224, 4.324907, 4.342075, 
    4.335614, 4.347477, 4.349862, 4.331839, 4.342902, 4.307461, 4.313179, 
    4.309772, 4.297355, 4.337106, 4.316681, 4.354437, 4.34334, 4.375771, 
    4.359628, 4.39137, 4.404985, 4.417808, 4.432834, 4.306675, 4.302355, 
    4.31009, 4.320809, 4.330761, 4.344017, 4.345373, 4.34786, 4.354303, 
    4.359725, 4.348649, 4.361084, 4.31451, 4.33888, 4.300725, 4.312197, 
    4.320176, 4.316672, 4.334875, 4.339172, 4.356662, 4.347614, 4.401625, 
    4.377684, 4.444284, 4.425619, 4.300847, 4.306659, 4.326927, 4.317276, 
    4.344901, 4.351717, 4.357261, 4.364357, 4.365122, 4.369329, 4.362436, 
    4.369056, 4.344045, 4.355212, 4.324604, 4.332044, 4.328619, 4.324867, 
    4.336455, 4.348824, 4.349084, 4.353055, 4.364265, 4.345013, 4.404728, 
    4.367803, 4.313002, 4.324226, 4.325825, 4.321476, 4.351034, 4.340311, 
    4.369226, 4.3614, 4.374227, 4.36785, 4.366913, 4.358732, 4.353644, 
    4.340803, 4.33037, 4.322105, 4.324026, 4.333107, 4.34958, 4.365193, 
    4.361771, 4.373251, 4.342895, 4.355611, 4.350695, 4.36352, 4.335443, 
    4.359358, 4.329344, 4.33197, 4.340098, 4.356478, 4.3601, 4.363976, 
    4.361583, 4.349998, 4.3481, 4.3399, 4.337639, 4.331398, 4.326236, 
    4.330953, 4.33591, 4.350001, 4.362724, 4.376617, 4.38002, 4.396302, 
    4.38305, 4.404935, 4.386334, 4.418557, 4.36074, 4.385779, 4.340467, 
    4.345335, 4.354152, 4.374403, 4.363459, 4.376257, 4.348025, 4.333423, 
    4.329645, 4.322608, 4.329806, 4.32922, 4.336113, 4.333897, 4.35047, 
    4.341563, 4.36689, 4.376155, 4.402372, 4.41849, 4.434923, 4.44219, 
    4.444403, 4.445329,
  3.964993, 3.978386, 3.975823, 3.986464, 3.980557, 3.98753, 3.967747, 
    3.978911, 3.971862, 3.966214, 4.007178, 3.986939, 4.02827, 4.015305, 
    4.047928, 4.026252, 4.052309, 4.047299, 4.062385, 4.058058, 4.077405, 
    4.064382, 4.087456, 4.074291, 4.076349, 4.063954, 3.991003, 4.004655, 
    3.990196, 3.99214, 3.991267, 3.98068, 3.975355, 3.963953, 3.96604, 
    3.974417, 3.993015, 3.986692, 4.002635, 4.002274, 4.020078, 4.012043, 
    4.042054, 4.033506, 4.058239, 4.052009, 4.057947, 4.056145, 4.05797, 
    4.048836, 4.052748, 4.044716, 4.013548, 4.02269, 3.99547, 3.979172, 
    3.968246, 3.960342, 3.961459, 3.963589, 3.974465, 3.984453, 3.992078, 
    3.997185, 4.002222, 4.017503, 4.025602, 4.043785, 4.040496, 4.046067, 
    4.051389, 4.060341, 4.058867, 4.062814, 4.045918, 4.057142, 4.038625, 
    4.043684, 4.003602, 3.988397, 3.981955, 3.976316, 3.962318, 3.972078, 
    3.968229, 3.977219, 3.982863, 3.980071, 3.997325, 3.990611, 4.026083, 
    4.010775, 4.050768, 4.041171, 4.053071, 4.046995, 4.05741, 4.048036, 
    4.064283, 4.067829, 4.065406, 4.074716, 4.047517, 4.057948, 3.979993, 
    3.980448, 3.982569, 3.973252, 3.972682, 3.963896, 3.971731, 3.974975, 
    3.98319, 3.988056, 3.992686, 4.002879, 4.014287, 4.030278, 4.041793, 
    4.049526, 4.044782, 4.04897, 4.044289, 4.042096, 4.066501, 4.052785, 
    4.073376, 4.072234, 4.062909, 4.072362, 3.980768, 3.978148, 3.968966, 
    3.976172, 3.962938, 3.970419, 3.97464, 3.990753, 3.994298, 3.997589, 
    4.004094, 4.012455, 4.027152, 4.039972, 4.051699, 4.050838, 4.051141, 
    4.053765, 4.047269, 4.054832, 4.056104, 4.052782, 4.072081, 4.06656, 
    4.07221, 4.068614, 3.978999, 3.983408, 3.981025, 3.985508, 3.98235, 
    3.996408, 4.00063, 4.020426, 4.01229, 4.025241, 4.013604, 4.015665, 
    4.025668, 4.014231, 4.039266, 4.022284, 4.053867, 4.036868, 4.054935, 
    4.051648, 4.05709, 4.061969, 4.068111, 4.079466, 4.076835, 4.086342, 
    3.989988, 3.995721, 3.995214, 4.001217, 4.005662, 4.015307, 4.030813, 
    4.024976, 4.035694, 4.037849, 4.021566, 4.03156, 3.999559, 4.004718, 
    4.001645, 3.990441, 4.026323, 4.00788, 4.041984, 4.031956, 4.061273, 
    4.046676, 4.075387, 4.087711, 4.099326, 4.11294, 3.99885, 3.994952, 
    4.001931, 4.011606, 4.020593, 4.032567, 4.033792, 4.03604, 4.041862, 
    4.046764, 4.036752, 4.047993, 4.005919, 4.027926, 3.99348, 4.003832, 
    4.011035, 4.007872, 4.024309, 4.028191, 4.043994, 4.035818, 4.084669, 
    4.063003, 4.123322, 4.106401, 3.993591, 3.998835, 4.01713, 4.008418, 
    4.033366, 4.039526, 4.044537, 4.050951, 4.051643, 4.055448, 4.049215, 
    4.055201, 4.032592, 4.042684, 4.015034, 4.021751, 4.01866, 4.015271, 
    4.025736, 4.03691, 4.037146, 4.040735, 4.050865, 4.033467, 4.087477, 
    4.054065, 4.00456, 4.014691, 4.016136, 4.012208, 4.038908, 4.029219, 
    4.055355, 4.048278, 4.059876, 4.05411, 4.053263, 4.045866, 4.041267, 
    4.029664, 4.02024, 4.012778, 4.014512, 4.022712, 4.037594, 4.051707, 
    4.048613, 4.058994, 4.031553, 4.043045, 4.038601, 4.050194, 4.024822, 
    4.04643, 4.019313, 4.021685, 4.029027, 4.043827, 4.047102, 4.050607, 
    4.048444, 4.037971, 4.036256, 4.028848, 4.026805, 4.021168, 4.016507, 
    4.020766, 4.025244, 4.037975, 4.049475, 4.062039, 4.065117, 4.079849, 
    4.067858, 4.087664, 4.070827, 4.100002, 4.04768, 4.070326, 4.02936, 
    4.033758, 4.041725, 4.060035, 4.050139, 4.061713, 4.036189, 4.022997, 
    4.019585, 4.013232, 4.019731, 4.019202, 4.025427, 4.023426, 4.038398, 
    4.03035, 4.053242, 4.06162, 4.085346, 4.099943, 4.114835, 4.121423, 
    4.12343, 4.124269,
  3.777921, 3.791298, 3.788693, 3.799511, 3.793505, 3.800595, 3.780629, 
    3.791831, 3.784675, 3.779123, 3.820599, 3.799994, 3.841569, 3.82876, 
    3.861022, 3.839573, 3.865362, 3.860399, 3.875352, 3.871062, 3.89026, 
    3.877334, 3.900249, 3.887167, 3.889211, 3.876908, 3.80413, 3.818028, 
    3.803308, 3.805286, 3.804398, 3.79363, 3.788217, 3.7769, 3.778951, 
    3.787264, 3.806176, 3.799744, 3.815973, 3.815605, 3.833474, 3.82554, 
    3.855206, 3.846749, 3.871241, 3.865066, 3.870951, 3.869165, 3.870974, 
    3.861922, 3.865798, 3.857842, 3.827025, 3.836055, 3.808676, 3.792095, 
    3.78112, 3.773352, 3.774449, 3.776542, 3.787313, 3.797467, 3.805224, 
    3.810423, 3.815552, 3.830929, 3.838932, 3.856919, 3.853665, 3.859179, 
    3.864452, 3.873325, 3.871863, 3.875778, 3.859032, 3.870153, 3.851813, 
    3.85682, 3.816955, 3.801478, 3.794925, 3.789194, 3.775293, 3.784888, 
    3.781102, 3.790112, 3.79585, 3.793011, 3.810565, 3.803731, 3.839406, 
    3.824268, 3.863837, 3.854332, 3.866118, 3.860099, 3.870419, 3.86113, 
    3.877235, 3.880753, 3.878349, 3.88759, 3.860615, 3.870951, 3.792932, 
    3.793394, 3.795551, 3.786081, 3.785502, 3.776844, 3.784546, 3.787831, 
    3.796182, 3.801132, 3.805843, 3.816222, 3.827755, 3.843554, 3.854948, 
    3.862606, 3.857908, 3.862055, 3.857419, 3.855248, 3.879435, 3.865834, 
    3.886259, 3.885126, 3.875871, 3.885253, 3.793719, 3.791056, 3.781827, 
    3.789048, 3.775902, 3.783256, 3.787491, 3.803875, 3.807483, 3.810834, 
    3.817459, 3.825946, 3.840465, 3.853145, 3.864758, 3.863906, 3.864206, 
    3.866806, 3.86037, 3.867864, 3.869124, 3.865832, 3.884974, 3.879495, 
    3.885102, 3.881533, 3.791922, 3.796404, 3.793982, 3.798539, 3.795328, 
    3.80963, 3.813929, 3.833817, 3.825783, 3.838575, 3.82708, 3.829115, 
    3.838996, 3.8277, 3.852446, 3.835653, 3.866907, 3.850072, 3.867965, 
    3.864708, 3.870101, 3.874939, 3.881034, 3.892308, 3.889694, 3.899142, 
    3.803097, 3.808931, 3.808416, 3.814529, 3.819057, 3.828762, 3.844084, 
    3.838314, 3.848912, 3.851044, 3.834945, 3.844822, 3.81284, 3.818094, 
    3.814964, 3.803558, 3.839645, 3.821316, 3.855137, 3.845214, 3.874249, 
    3.859782, 3.888256, 3.900501, 3.912058, 3.925619, 3.812118, 3.808149, 
    3.815257, 3.825108, 3.833983, 3.845819, 3.847031, 3.849254, 3.855017, 
    3.85987, 3.849958, 3.861087, 3.819317, 3.841229, 3.806651, 3.817192, 
    3.824533, 3.821309, 3.837655, 3.841492, 3.857127, 3.849035, 3.897476, 
    3.875964, 3.935974, 3.919103, 3.806764, 3.812103, 3.830562, 3.821865, 
    3.84661, 3.852704, 3.857664, 3.864017, 3.864703, 3.868473, 3.862298, 
    3.868229, 3.845844, 3.85583, 3.828492, 3.835128, 3.832073, 3.828727, 
    3.839065, 3.850115, 3.850349, 3.8539, 3.863929, 3.84671, 3.900266, 
    3.8671, 3.817935, 3.828153, 3.82958, 3.825703, 3.852093, 3.842508, 
    3.868381, 3.86137, 3.872864, 3.867148, 3.866308, 3.858981, 3.854427, 
    3.842948, 3.833634, 3.826265, 3.827977, 3.836076, 3.850791, 3.864766, 
    3.861701, 3.871989, 3.844817, 3.856187, 3.851789, 3.863268, 3.838161, 
    3.859536, 3.832719, 3.835062, 3.842318, 3.856961, 3.860205, 3.863677, 
    3.861534, 3.851165, 3.849468, 3.842141, 3.840122, 3.834552, 3.829947, 
    3.834154, 3.838578, 3.851169, 3.862554, 3.875009, 3.878062, 3.892686, 
    3.88078, 3.900452, 3.883724, 3.912728, 3.860775, 3.88323, 3.842648, 
    3.846997, 3.85488, 3.87302, 3.863214, 3.874684, 3.849402, 3.836357, 
    3.832988, 3.826713, 3.833131, 3.832609, 3.83876, 3.836782, 3.851588, 
    3.843627, 3.866287, 3.874593, 3.898151, 3.912671, 3.927509, 3.93408, 
    3.936082, 3.93692,
  3.838243, 3.85263, 3.849826, 3.861443, 3.855007, 3.862575, 3.841152, 
    3.853203, 3.845504, 3.839534, 3.883493, 3.861948, 3.906065, 3.892179, 
    3.927207, 3.9039, 3.931933, 3.92653, 3.942823, 3.938144, 3.959105, 
    3.944985, 3.970038, 3.955725, 3.957959, 3.944521, 3.866267, 3.880801, 
    3.865409, 3.867476, 3.866548, 3.855141, 3.849313, 3.837145, 3.83935, 
    3.848288, 3.868405, 3.861687, 3.878651, 3.878266, 3.897287, 3.888693, 
    3.92088, 3.911689, 3.938339, 3.93161, 3.938023, 3.936077, 3.938048, 
    3.928187, 3.932407, 3.923747, 3.890301, 3.900084, 3.871018, 3.853488, 
    3.84168, 3.833335, 3.834513, 3.836761, 3.848341, 3.859274, 3.867411, 
    3.872845, 3.878211, 3.894528, 3.903204, 3.922743, 3.919204, 3.925201, 
    3.930942, 3.940612, 3.939017, 3.943287, 3.925041, 3.937153, 3.917191, 
    3.922635, 3.879677, 3.863497, 3.856535, 3.850365, 3.835419, 3.845732, 
    3.841662, 3.851354, 3.857532, 3.854474, 3.872994, 3.86585, 3.903719, 
    3.887337, 3.930271, 3.91993, 3.932756, 3.926203, 3.937443, 3.927325, 
    3.944878, 3.948717, 3.946093, 3.956187, 3.926765, 3.938024, 3.854389, 
    3.854887, 3.85721, 3.847015, 3.846392, 3.837085, 3.845365, 3.848899, 
    3.85789, 3.863136, 3.868057, 3.878911, 3.891091, 3.90822, 3.920599, 
    3.928931, 3.923818, 3.928332, 3.923287, 3.920926, 3.947278, 3.932447, 
    3.954733, 3.953494, 3.943389, 3.953634, 3.855237, 3.85237, 3.842441, 
    3.850208, 3.836074, 3.843977, 3.848532, 3.866001, 3.869771, 3.873275, 
    3.880207, 3.889132, 3.904867, 3.918638, 3.931276, 3.930348, 3.930675, 
    3.933506, 3.926498, 3.934659, 3.936031, 3.932445, 3.953328, 3.947344, 
    3.953468, 3.949569, 3.853302, 3.85813, 3.85552, 3.860429, 3.85697, 
    3.872016, 3.876512, 3.897658, 3.888957, 3.902817, 3.890361, 3.892564, 
    3.903273, 3.891032, 3.917878, 3.899648, 3.933616, 3.915298, 3.934769, 
    3.931221, 3.937097, 3.942373, 3.949024, 3.961346, 3.958487, 3.968826, 
    3.865188, 3.871285, 3.870747, 3.87714, 3.88188, 3.892182, 3.908795, 
    3.902534, 3.914039, 3.916356, 3.898881, 3.909597, 3.875372, 3.880871, 
    3.877595, 3.865669, 3.903977, 3.884245, 3.920804, 3.910022, 3.94162, 
    3.925857, 3.956915, 3.970315, 3.982987, 3.997886, 3.874617, 3.870468, 
    3.877902, 3.888225, 3.897839, 3.910679, 3.911996, 3.91441, 3.920674, 
    3.925953, 3.915175, 3.927279, 3.88215, 3.905697, 3.868902, 3.879926, 
    3.887615, 3.884238, 3.90182, 3.905982, 3.922968, 3.914172, 3.967002, 
    3.94349, 4.009287, 3.990723, 3.86902, 3.874603, 3.894131, 3.88482, 
    3.911538, 3.918159, 3.923554, 3.930469, 3.931216, 3.935323, 3.928596, 
    3.935056, 3.910706, 3.921558, 3.89189, 3.899079, 3.895769, 3.892144, 
    3.903349, 3.915345, 3.9156, 3.91946, 3.93037, 3.911647, 3.970056, 
    3.933825, 3.880704, 3.891521, 3.893068, 3.88887, 3.917495, 3.907085, 
    3.935222, 3.927586, 3.94011, 3.933879, 3.932963, 3.924986, 3.920033, 
    3.907562, 3.89746, 3.889478, 3.891332, 3.900108, 3.91608, 3.931284, 
    3.927946, 3.939156, 3.909591, 3.921946, 3.917164, 3.929652, 3.902369, 
    3.925588, 3.896469, 3.899008, 3.906879, 3.922788, 3.926318, 3.930097, 
    3.927764, 3.916487, 3.914643, 3.906687, 3.904495, 3.898455, 3.893466, 
    3.898024, 3.902821, 3.916491, 3.928875, 3.942448, 3.94578, 3.961759, 
    3.948746, 3.970259, 3.951961, 3.983721, 3.926938, 3.951421, 3.907237, 
    3.911959, 3.920525, 3.940279, 3.929593, 3.942094, 3.914571, 3.900412, 
    3.89676, 3.889963, 3.896915, 3.896349, 3.903018, 3.900873, 3.916946, 
    3.908299, 3.932941, 3.941995, 3.967741, 3.983659, 3.999966, 4.007201, 
    4.009407, 4.01033,
  3.964783, 3.983002, 3.979445, 3.994249, 3.986021, 3.995738, 3.968461, 
    3.98373, 3.973967, 3.966415, 4.023345, 3.994913, 4.052799, 4.034864, 
    4.080283, 4.049997, 4.086456, 4.0794, 4.100724, 4.094587, 4.122168, 
    4.103564, 4.136643, 4.117705, 4.120654, 4.102954, 4.000596, 4.01978, 
    3.999466, 4.002187, 4.000965, 3.986191, 3.978794, 3.963398, 3.966182, 
    3.977495, 4.003412, 3.99457, 4.016936, 4.016428, 4.041451, 4.03024, 
    4.072035, 4.060089, 4.094842, 4.086035, 4.094428, 4.091878, 4.094461, 
    4.081562, 4.087077, 4.07577, 4.032374, 4.045063, 4.006856, 3.984092, 
    3.969128, 3.958588, 3.960075, 3.962912, 3.977561, 3.991446, 4.002102, 
    4.009266, 4.016355, 4.037891, 4.049096, 4.074462, 4.069854, 4.077666, 
    4.085161, 4.097823, 4.095732, 4.101334, 4.077458, 4.093288, 4.067235, 
    4.074321, 4.018293, 3.99695, 3.987963, 3.980129, 3.961218, 3.974256, 
    3.969105, 3.981383, 3.98923, 3.985344, 4.009463, 4.000047, 4.049763, 
    4.028441, 4.084285, 4.070798, 4.087533, 4.078973, 4.093668, 4.080437, 
    4.103423, 4.108471, 4.10502, 4.118315, 4.079706, 4.094429, 3.985236, 
    3.985869, 3.988821, 3.975882, 3.975093, 3.963321, 3.973791, 3.978269, 
    3.989686, 3.996475, 4.002953, 4.017281, 4.033423, 4.055591, 4.07167, 
    4.082534, 4.075863, 4.081752, 4.075171, 4.072095, 4.106578, 4.087129, 
    4.116396, 4.114763, 4.101468, 4.114947, 3.986314, 3.982672, 3.970091, 
    3.979929, 3.962044, 3.972034, 3.977804, 4.000245, 4.005212, 4.009833, 
    4.018994, 4.030823, 4.051249, 4.069118, 4.085598, 4.084384, 4.084812, 
    4.088514, 4.079359, 4.090022, 4.091819, 4.087126, 4.114544, 4.106665, 
    4.114728, 4.109593, 3.983855, 3.98999, 3.986672, 3.992917, 3.988516, 
    4.008172, 4.014109, 4.04193, 4.03059, 4.048596, 4.032454, 4.03536, 
    4.049186, 4.033345, 4.068129, 4.044499, 4.088658, 4.064775, 4.090167, 
    4.085526, 4.093215, 4.100133, 4.108875, 4.12513, 4.121352, 4.135036, 
    3.999175, 4.007208, 4.006498, 4.014939, 4.021208, 4.034868, 4.056336, 
    4.048231, 4.06314, 4.06615, 4.04351, 4.057375, 4.012603, 4.019874, 
    4.01554, 3.999808, 4.050097, 4.024341, 4.071937, 4.057928, 4.099145, 
    4.078522, 4.119276, 4.13701, 4.153869, 4.173799, 4.011606, 4.00613, 
    4.015945, 4.029619, 4.042163, 4.058779, 4.060488, 4.063622, 4.071768, 
    4.078648, 4.064616, 4.080377, 4.021566, 4.052323, 4.004066, 4.018622, 
    4.028809, 4.024332, 4.047307, 4.052692, 4.074756, 4.063313, 4.132617, 
    4.1016, 4.189131, 4.164202, 4.004221, 4.011586, 4.03738, 4.025104, 
    4.059893, 4.068495, 4.075519, 4.084542, 4.085519, 4.090891, 4.082097, 
    4.090542, 4.058815, 4.072919, 4.034485, 4.043765, 4.039493, 4.034819, 
    4.049285, 4.064836, 4.065168, 4.070187, 4.084414, 4.060035, 4.136666, 
    4.088931, 4.019652, 4.033996, 4.03601, 4.030475, 4.067631, 4.054121, 
    4.09076, 4.080778, 4.097164, 4.089002, 4.087804, 4.077385, 4.070932, 
    4.054738, 4.041675, 4.031282, 4.033744, 4.045094, 4.065792, 4.085608, 
    4.081247, 4.095913, 4.057368, 4.073424, 4.067201, 4.083476, 4.048017, 
    4.078171, 4.040396, 4.043674, 4.053854, 4.07452, 4.079124, 4.084057, 
    4.081011, 4.06632, 4.063924, 4.053605, 4.050767, 4.042959, 4.036523, 
    4.042403, 4.048601, 4.066325, 4.082461, 4.100232, 4.104609, 4.125676, 
    4.10851, 4.136936, 4.112742, 4.154847, 4.079932, 4.112031, 4.054317, 
    4.06044, 4.071573, 4.097386, 4.083399, 4.099767, 4.06383, 4.045487, 
    4.040771, 4.031926, 4.040972, 4.040241, 4.048857, 4.046083, 4.066917, 
    4.055694, 4.087775, 4.099637, 4.133597, 4.154765, 4.176591, 4.18632, 
    4.189293, 4.190537,
  4.394931, 4.425735, 4.419685, 4.444981, 4.430883, 4.447541, 4.401113, 
    4.426975, 4.410401, 4.397671, 4.495613, 4.446121, 4.549213, 4.516021, 
    4.601168, 4.543991, 4.612795, 4.599476, 4.639682, 4.628071, 4.680817, 
    4.64508, 4.709098, 4.672182, 4.677884, 4.643919, 4.455919, 4.489343, 
    4.453968, 4.458671, 4.456557, 4.431174, 4.41858, 4.392606, 4.39728, 
    4.416376, 4.460792, 4.445531, 4.484354, 4.483463, 4.528148, 4.507799, 
    4.585434, 4.562863, 4.628553, 4.612007, 4.627772, 4.622969, 4.627834, 
    4.60362, 4.613957, 4.592544, 4.511585, 4.53483, 4.466766, 4.427591, 
    4.402236, 4.384558, 4.387042, 4.391791, 4.416488, 4.440166, 4.458524, 
    4.470959, 4.483335, 4.521585, 4.542316, 4.590051, 4.581295, 4.596162, 
    4.610373, 4.634184, 4.630231, 4.64084, 4.595766, 4.625624, 4.576335, 
    4.589783, 4.486733, 4.449629, 4.434201, 4.420846, 4.388955, 4.41089, 
    4.402197, 4.422978, 4.436369, 4.429728, 4.471301, 4.454971, 4.543556, 
    4.504612, 4.608737, 4.583086, 4.614812, 4.59866, 4.626339, 4.601462, 
    4.644811, 4.654441, 4.647852, 4.67336, 4.600064, 4.627773, 4.429543, 
    4.430624, 4.435669, 4.413641, 4.412306, 4.392478, 4.410104, 4.417688, 
    4.43715, 4.44881, 4.459997, 4.484957, 4.51345, 4.554431, 4.58474, 
    4.605471, 4.592722, 4.603983, 4.591402, 4.585548, 4.650825, 4.614055, 
    4.669657, 4.666512, 4.641094, 4.666865, 4.431383, 4.425173, 4.403858, 
    4.420507, 4.390338, 4.407135, 4.4169, 4.455313, 4.463913, 4.471945, 
    4.487963, 4.508832, 4.546323, 4.579899, 4.61119, 4.608923, 4.60972, 
    4.616651, 4.599398, 4.61948, 4.622858, 4.614048, 4.666091, 4.65099, 
    4.666445, 4.656587, 4.427188, 4.437671, 4.431995, 4.44269, 4.435147, 
    4.469054, 4.479405, 4.529032, 4.508419, 4.541387, 4.511726, 4.516931, 
    4.542483, 4.51331, 4.578026, 4.533785, 4.616921, 4.571688, 4.619751, 
    4.611056, 4.625486, 4.638561, 4.655214, 4.68657, 4.679235, 4.705936, 
    4.453466, 4.467378, 4.466145, 4.480857, 4.491853, 4.516028, 4.555826, 
    4.540708, 4.568604, 4.574283, 4.531953, 4.557772, 4.476775, 4.489507, 
    4.481909, 4.454559, 4.544178, 4.49737, 4.585248, 4.558807, 4.636688, 
    4.597797, 4.675217, 4.70982, 4.743316, 4.783701, 4.475035, 4.465506, 
    4.482618, 4.506698, 4.529464, 4.560404, 4.563612, 4.569513, 4.584926, 
    4.598038, 4.571386, 4.601347, 4.492483, 4.548326, 4.461925, 4.487311, 
    4.505264, 4.497354, 4.538991, 4.549014, 4.590611, 4.56893, 4.701188, 
    4.641345, 4.815381, 4.764145, 4.462195, 4.475001, 4.520644, 4.498715, 
    4.562496, 4.578719, 4.592064, 4.609218, 4.611042, 4.621113, 4.604644, 
    4.620458, 4.560471, 4.587114, 4.515338, 4.532426, 4.524535, 4.515938, 
    4.542666, 4.571802, 4.572429, 4.581925, 4.608977, 4.562761, 4.709143, 
    4.617431, 4.489119, 4.514466, 4.518125, 4.508215, 4.577083, 4.551681, 
    4.620866, 4.602116, 4.632938, 4.617564, 4.615319, 4.595627, 4.58334, 
    4.552835, 4.528562, 4.509647, 4.514019, 4.534887, 4.573606, 4.611209, 
    4.603016, 4.630574, 4.557758, 4.588075, 4.57627, 4.607226, 4.540309, 
    4.597127, 4.5262, 4.532257, 4.551182, 4.590161, 4.598949, 4.608312, 
    4.602562, 4.574605, 4.570083, 4.550718, 4.545427, 4.530935, 4.519067, 
    4.529907, 4.541395, 4.574615, 4.605334, 4.638749, 4.647069, 4.687633, 
    4.654514, 4.709675, 4.662626, 4.745277, 4.600495, 4.661262, 4.552049, 
    4.563523, 4.584557, 4.633358, 4.607083, 4.637867, 4.569905, 4.535615, 
    4.526893, 4.51079, 4.527263, 4.525915, 4.541871, 4.53672, 4.575733, 
    4.554623, 4.615264, 4.63762, 4.703111, 4.745113, 4.789431, 4.809532, 
    4.815718, 4.818313,
  6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465,
  6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  25080.91, 25097.15, 25093.97, 25107.23, 25099.85, 25108.56, 25084.18, 
    25097.8, 25089.09, 25082.36, 25133.43, 25107.82, 25160.68, 25143.89, 
    25186.69, 25158.05, 25192.51, 25185.85, 25205.97, 25200.17, 25226.39, 
    25208.66, 25240.3, 25222.12, 25224.94, 25208.08, 25112.92, 25130.21, 
    25111.9, 25114.35, 25113.25, 25100.01, 25093.39, 25079.68, 25082.15, 
    25092.23, 25115.45, 25107.51, 25127.63, 25127.17, 25150.04, 25139.69, 
    25178.85, 25167.54, 25200.41, 25192.12, 25200.02, 25197.62, 25200.05, 
    25187.91, 25193.1, 25182.39, 25141.62, 25153.42, 25118.54, 25098.13, 
    25084.78, 25075.41, 25076.73, 25079.25, 25092.29, 25104.71, 25114.27, 
    25120.71, 25127.11, 25146.72, 25157.2, 25181.15, 25176.78, 25184.2, 
    25191.29, 25203.23, 25201.25, 25206.55, 25184, 25198.95, 25174.3, 
    25181.02, 25128.86, 25109.65, 25101.59, 25094.58, 25077.74, 25089.35, 
    25084.75, 25095.71, 25102.73, 25099.25, 25120.89, 25112.42, 25157.83, 
    25138.05, 25190.47, 25177.67, 25193.52, 25185.44, 25199.3, 25186.83, 
    25208.53, 25213.32, 25210.04, 25222.7, 25186.14, 25200.02, 25099.15, 
    25099.72, 25102.36, 25090.79, 25090.09, 25079.61, 25088.93, 25092.92, 
    25103.13, 25109.22, 25115.03, 25127.95, 25142.58, 25163.31, 25178.5, 
    25188.83, 25182.48, 25188.09, 25181.82, 25178.9, 25211.52, 25193.14, 
    25220.87, 25219.31, 25206.68, 25219.49, 25100.12, 25096.86, 25085.63, 
    25094.41, 25078.48, 25087.36, 25092.51, 25112.6, 25117.06, 25121.22, 
    25129.49, 25140.22, 25159.22, 25176.08, 25191.71, 25190.56, 25190.97, 
    25194.45, 25185.81, 25195.87, 25197.56, 25193.14, 25219.1, 25211.6, 
    25219.28, 25214.39, 25097.91, 25103.41, 25100.44, 25106.03, 25102.09, 
    25119.73, 25125.08, 25150.49, 25140.01, 25156.73, 25141.7, 25144.35, 
    25157.29, 25142.51, 25175.14, 25152.89, 25194.58, 25171.97, 25196, 
    25191.64, 25198.88, 25205.41, 25213.71, 25229.22, 25225.61, 25238.75, 
    25111.64, 25118.86, 25118.22, 25125.83, 25131.5, 25143.89, 25164.01, 
    25156.39, 25170.43, 25173.27, 25151.97, 25164.99, 25123.72, 25130.29, 
    25126.37, 25112.21, 25158.14, 25134.34, 25178.75, 25165.51, 25204.48, 
    25185.01, 25223.62, 25240.65, 25257.01, 25276.54, 25122.82, 25117.89, 
    25126.74, 25139.12, 25150.71, 25166.31, 25167.92, 25170.88, 25178.59, 
    25185.13, 25171.82, 25186.78, 25131.82, 25160.23, 25116.03, 25129.16, 
    25138.39, 25134.33, 25155.53, 25160.58, 25181.43, 25170.59, 25236.42, 
    25206.8, 25291.73, 25267.11, 25116.17, 25122.8, 25146.24, 25135.03, 
    25167.36, 25175.49, 25182.15, 25190.71, 25191.63, 25196.69, 25188.41, 
    25196.36, 25166.34, 25179.69, 25143.54, 25152.21, 25148.21, 25143.85, 
    25157.38, 25172.03, 25172.34, 25177.09, 25190.59, 25167.49, 25240.32, 
    25194.84, 25130.09, 25143.1, 25144.96, 25139.9, 25174.67, 25161.92, 
    25196.56, 25187.16, 25202.6, 25194.91, 25193.78, 25183.93, 25177.8, 
    25162.51, 25150.25, 25140.63, 25142.87, 25153.45, 25172.93, 25191.71, 
    25187.61, 25201.42, 25164.98, 25180.16, 25174.27, 25189.71, 25156.19, 
    25184.68, 25149.05, 25152.12, 25161.67, 25181.21, 25185.58, 25190.26, 
    25187.38, 25173.43, 25171.17, 25161.44, 25158.77, 25151.45, 25145.44, 
    25150.93, 25156.74, 25173.44, 25188.76, 25205.51, 25209.65, 25229.75, 
    25213.36, 25240.58, 25217.38, 25257.96, 25186.35, 25216.71, 25162.11, 
    25167.88, 25178.41, 25202.81, 25189.64, 25205.07, 25171.08, 25153.82, 
    25149.41, 25141.22, 25149.59, 25148.91, 25156.98, 25154.38, 25174, 
    25163.4, 25193.75, 25204.94, 25237.36, 25257.88, 25279.3, 25288.94, 
    25291.89, 25293.13 ;

 HCSOI =
  25080.91, 25097.15, 25093.97, 25107.23, 25099.85, 25108.56, 25084.18, 
    25097.8, 25089.09, 25082.36, 25133.43, 25107.82, 25160.68, 25143.89, 
    25186.69, 25158.05, 25192.51, 25185.85, 25205.97, 25200.17, 25226.39, 
    25208.66, 25240.3, 25222.12, 25224.94, 25208.08, 25112.92, 25130.21, 
    25111.9, 25114.35, 25113.25, 25100.01, 25093.39, 25079.68, 25082.15, 
    25092.23, 25115.45, 25107.51, 25127.63, 25127.17, 25150.04, 25139.69, 
    25178.85, 25167.54, 25200.41, 25192.12, 25200.02, 25197.62, 25200.05, 
    25187.91, 25193.1, 25182.39, 25141.62, 25153.42, 25118.54, 25098.13, 
    25084.78, 25075.41, 25076.73, 25079.25, 25092.29, 25104.71, 25114.27, 
    25120.71, 25127.11, 25146.72, 25157.2, 25181.15, 25176.78, 25184.2, 
    25191.29, 25203.23, 25201.25, 25206.55, 25184, 25198.95, 25174.3, 
    25181.02, 25128.86, 25109.65, 25101.59, 25094.58, 25077.74, 25089.35, 
    25084.75, 25095.71, 25102.73, 25099.25, 25120.89, 25112.42, 25157.83, 
    25138.05, 25190.47, 25177.67, 25193.52, 25185.44, 25199.3, 25186.83, 
    25208.53, 25213.32, 25210.04, 25222.7, 25186.14, 25200.02, 25099.15, 
    25099.72, 25102.36, 25090.79, 25090.09, 25079.61, 25088.93, 25092.92, 
    25103.13, 25109.22, 25115.03, 25127.95, 25142.58, 25163.31, 25178.5, 
    25188.83, 25182.48, 25188.09, 25181.82, 25178.9, 25211.52, 25193.14, 
    25220.87, 25219.31, 25206.68, 25219.49, 25100.12, 25096.86, 25085.63, 
    25094.41, 25078.48, 25087.36, 25092.51, 25112.6, 25117.06, 25121.22, 
    25129.49, 25140.22, 25159.22, 25176.08, 25191.71, 25190.56, 25190.97, 
    25194.45, 25185.81, 25195.87, 25197.56, 25193.14, 25219.1, 25211.6, 
    25219.28, 25214.39, 25097.91, 25103.41, 25100.44, 25106.03, 25102.09, 
    25119.73, 25125.08, 25150.49, 25140.01, 25156.73, 25141.7, 25144.35, 
    25157.29, 25142.51, 25175.14, 25152.89, 25194.58, 25171.97, 25196, 
    25191.64, 25198.88, 25205.41, 25213.71, 25229.22, 25225.61, 25238.75, 
    25111.64, 25118.86, 25118.22, 25125.83, 25131.5, 25143.89, 25164.01, 
    25156.39, 25170.43, 25173.27, 25151.97, 25164.99, 25123.72, 25130.29, 
    25126.37, 25112.21, 25158.14, 25134.34, 25178.75, 25165.51, 25204.48, 
    25185.01, 25223.62, 25240.65, 25257.01, 25276.54, 25122.82, 25117.89, 
    25126.74, 25139.12, 25150.71, 25166.31, 25167.92, 25170.88, 25178.59, 
    25185.13, 25171.82, 25186.78, 25131.82, 25160.23, 25116.03, 25129.16, 
    25138.39, 25134.33, 25155.53, 25160.58, 25181.43, 25170.59, 25236.42, 
    25206.8, 25291.73, 25267.11, 25116.17, 25122.8, 25146.24, 25135.03, 
    25167.36, 25175.49, 25182.15, 25190.71, 25191.63, 25196.69, 25188.41, 
    25196.36, 25166.34, 25179.69, 25143.54, 25152.21, 25148.21, 25143.85, 
    25157.38, 25172.03, 25172.34, 25177.09, 25190.59, 25167.49, 25240.32, 
    25194.84, 25130.09, 25143.1, 25144.96, 25139.9, 25174.67, 25161.92, 
    25196.56, 25187.16, 25202.6, 25194.91, 25193.78, 25183.93, 25177.8, 
    25162.51, 25150.25, 25140.63, 25142.87, 25153.45, 25172.93, 25191.71, 
    25187.61, 25201.42, 25164.98, 25180.16, 25174.27, 25189.71, 25156.19, 
    25184.68, 25149.05, 25152.12, 25161.67, 25181.21, 25185.58, 25190.26, 
    25187.38, 25173.43, 25171.17, 25161.44, 25158.77, 25151.45, 25145.44, 
    25150.93, 25156.74, 25173.44, 25188.76, 25205.51, 25209.65, 25229.75, 
    25213.36, 25240.58, 25217.38, 25257.96, 25186.35, 25216.71, 25162.11, 
    25167.88, 25178.41, 25202.81, 25189.64, 25205.07, 25171.08, 25153.82, 
    25149.41, 25141.22, 25149.59, 25148.91, 25156.98, 25154.38, 25174, 
    25163.4, 25193.75, 25204.94, 25237.36, 25257.88, 25279.3, 25288.94, 
    25291.89, 25293.13 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  7.623649e-08, 7.644516e-08, 7.640461e-08, 7.657286e-08, 7.647954e-08, 
    7.658971e-08, 7.627882e-08, 7.645342e-08, 7.634197e-08, 7.62553e-08, 
    7.689925e-08, 7.658038e-08, 7.723048e-08, 7.70272e-08, 7.753781e-08, 
    7.719884e-08, 7.760615e-08, 7.752807e-08, 7.776314e-08, 7.76958e-08, 
    7.799632e-08, 7.779421e-08, 7.815211e-08, 7.794808e-08, 7.797998e-08, 
    7.778754e-08, 7.664459e-08, 7.685954e-08, 7.663184e-08, 7.66625e-08, 
    7.664875e-08, 7.648146e-08, 7.639712e-08, 7.622056e-08, 7.625263e-08, 
    7.638231e-08, 7.667629e-08, 7.657653e-08, 7.682798e-08, 7.682231e-08, 
    7.710213e-08, 7.697598e-08, 7.744618e-08, 7.731258e-08, 7.769862e-08, 
    7.760154e-08, 7.769405e-08, 7.766601e-08, 7.769442e-08, 7.755205e-08, 
    7.761304e-08, 7.748777e-08, 7.69996e-08, 7.714308e-08, 7.671504e-08, 
    7.64575e-08, 7.628647e-08, 7.616506e-08, 7.618222e-08, 7.621494e-08, 
    7.638307e-08, 7.654115e-08, 7.666159e-08, 7.674213e-08, 7.682149e-08, 
    7.706157e-08, 7.718869e-08, 7.747317e-08, 7.742187e-08, 7.750881e-08, 
    7.759189e-08, 7.773131e-08, 7.770838e-08, 7.776979e-08, 7.750653e-08, 
    7.768149e-08, 7.739264e-08, 7.747165e-08, 7.684295e-08, 7.660345e-08, 
    7.650154e-08, 7.64124e-08, 7.619542e-08, 7.634526e-08, 7.628619e-08, 
    7.642673e-08, 7.651601e-08, 7.647186e-08, 7.674434e-08, 7.663841e-08, 
    7.719622e-08, 7.695601e-08, 7.758219e-08, 7.74324e-08, 7.76181e-08, 
    7.752336e-08, 7.768568e-08, 7.75396e-08, 7.779266e-08, 7.784774e-08, 
    7.781009e-08, 7.795472e-08, 7.753149e-08, 7.769404e-08, 7.647062e-08, 
    7.647782e-08, 7.651137e-08, 7.636387e-08, 7.635484e-08, 7.621968e-08, 
    7.633997e-08, 7.639117e-08, 7.65212e-08, 7.659807e-08, 7.667116e-08, 
    7.683181e-08, 7.701119e-08, 7.726197e-08, 7.744212e-08, 7.756284e-08, 
    7.748882e-08, 7.755416e-08, 7.748111e-08, 7.744688e-08, 7.782709e-08, 
    7.761361e-08, 7.793392e-08, 7.791621e-08, 7.777125e-08, 7.791819e-08, 
    7.648288e-08, 7.644144e-08, 7.629752e-08, 7.641015e-08, 7.620496e-08, 
    7.631981e-08, 7.638584e-08, 7.66406e-08, 7.669659e-08, 7.674847e-08, 
    7.685095e-08, 7.698243e-08, 7.721304e-08, 7.741363e-08, 7.759672e-08, 
    7.758331e-08, 7.758803e-08, 7.762892e-08, 7.752763e-08, 7.764555e-08, 
    7.766533e-08, 7.76136e-08, 7.791383e-08, 7.782807e-08, 7.791583e-08, 
    7.785999e-08, 7.645492e-08, 7.652464e-08, 7.648696e-08, 7.65578e-08, 
    7.650789e-08, 7.672979e-08, 7.679631e-08, 7.710752e-08, 7.697984e-08, 
    7.718307e-08, 7.700049e-08, 7.703284e-08, 7.718965e-08, 7.701037e-08, 
    7.740255e-08, 7.713665e-08, 7.76305e-08, 7.736501e-08, 7.764714e-08, 
    7.759594e-08, 7.768072e-08, 7.775665e-08, 7.785217e-08, 7.802836e-08, 
    7.798757e-08, 7.813491e-08, 7.662858e-08, 7.671898e-08, 7.671105e-08, 
    7.680566e-08, 7.687562e-08, 7.702726e-08, 7.727039e-08, 7.717897e-08, 
    7.73468e-08, 7.738048e-08, 7.712552e-08, 7.728205e-08, 7.67795e-08, 
    7.686069e-08, 7.681236e-08, 7.66357e-08, 7.720001e-08, 7.691045e-08, 
    7.744509e-08, 7.728828e-08, 7.774582e-08, 7.751829e-08, 7.796511e-08, 
    7.815598e-08, 7.833569e-08, 7.854553e-08, 7.676834e-08, 7.670692e-08, 
    7.681692e-08, 7.696904e-08, 7.711023e-08, 7.729785e-08, 7.731705e-08, 
    7.735219e-08, 7.744323e-08, 7.751974e-08, 7.736328e-08, 7.753892e-08, 
    7.687949e-08, 7.722515e-08, 7.668368e-08, 7.684673e-08, 7.696008e-08, 
    7.691038e-08, 7.716854e-08, 7.722935e-08, 7.747646e-08, 7.734874e-08, 
    7.810886e-08, 7.777265e-08, 7.870533e-08, 7.844478e-08, 7.668545e-08, 
    7.676814e-08, 7.705584e-08, 7.691897e-08, 7.731038e-08, 7.740669e-08, 
    7.748498e-08, 7.758503e-08, 7.759585e-08, 7.765512e-08, 7.755798e-08, 
    7.765129e-08, 7.729825e-08, 7.745604e-08, 7.702298e-08, 7.71284e-08, 
    7.707991e-08, 7.702671e-08, 7.71909e-08, 7.736573e-08, 7.736951e-08, 
    7.742555e-08, 7.758342e-08, 7.731197e-08, 7.815218e-08, 7.763335e-08, 
    7.68583e-08, 7.701748e-08, 7.704026e-08, 7.697859e-08, 7.739703e-08, 
    7.724544e-08, 7.765367e-08, 7.754338e-08, 7.77241e-08, 7.76343e-08, 
    7.762108e-08, 7.750573e-08, 7.74339e-08, 7.725239e-08, 7.710467e-08, 
    7.698755e-08, 7.701478e-08, 7.714345e-08, 7.737644e-08, 7.759681e-08, 
    7.754854e-08, 7.771037e-08, 7.728201e-08, 7.746164e-08, 7.739221e-08, 
    7.757325e-08, 7.717654e-08, 7.751427e-08, 7.709018e-08, 7.712737e-08, 
    7.724243e-08, 7.74738e-08, 7.752503e-08, 7.757966e-08, 7.754596e-08, 
    7.738236e-08, 7.735557e-08, 7.723964e-08, 7.720762e-08, 7.711928e-08, 
    7.704612e-08, 7.711296e-08, 7.718313e-08, 7.738244e-08, 7.7562e-08, 
    7.775772e-08, 7.780563e-08, 7.803415e-08, 7.784809e-08, 7.815506e-08, 
    7.789401e-08, 7.834588e-08, 7.753389e-08, 7.788639e-08, 7.724768e-08, 
    7.731652e-08, 7.744099e-08, 7.772646e-08, 7.757239e-08, 7.775259e-08, 
    7.735452e-08, 7.714787e-08, 7.709443e-08, 7.699466e-08, 7.709671e-08, 
    7.708842e-08, 7.718606e-08, 7.715469e-08, 7.738906e-08, 7.726317e-08, 
    7.762075e-08, 7.775118e-08, 7.811946e-08, 7.834512e-08, 7.857481e-08, 
    7.867618e-08, 7.870703e-08, 7.871993e-08 ;

 HR_vr =
  2.780798e-07, 2.787892e-07, 2.786514e-07, 2.79223e-07, 2.789061e-07, 
    2.792802e-07, 2.782238e-07, 2.788173e-07, 2.784386e-07, 2.781439e-07, 
    2.803304e-07, 2.792485e-07, 2.814534e-07, 2.807647e-07, 2.824936e-07, 
    2.813461e-07, 2.827247e-07, 2.824608e-07, 2.832555e-07, 2.83028e-07, 
    2.840427e-07, 2.833605e-07, 2.845685e-07, 2.8388e-07, 2.839877e-07, 
    2.83338e-07, 2.794667e-07, 2.801957e-07, 2.794234e-07, 2.795274e-07, 
    2.794808e-07, 2.789126e-07, 2.786258e-07, 2.780257e-07, 2.781348e-07, 
    2.785756e-07, 2.795742e-07, 2.792356e-07, 2.800892e-07, 2.800699e-07, 
    2.810187e-07, 2.805911e-07, 2.821837e-07, 2.817316e-07, 2.830375e-07, 
    2.827093e-07, 2.83022e-07, 2.829273e-07, 2.830233e-07, 2.825419e-07, 
    2.827481e-07, 2.823245e-07, 2.806711e-07, 2.811574e-07, 2.797058e-07, 
    2.788309e-07, 2.782498e-07, 2.778369e-07, 2.778953e-07, 2.780066e-07, 
    2.785782e-07, 2.791154e-07, 2.795244e-07, 2.797978e-07, 2.800672e-07, 
    2.808809e-07, 2.813118e-07, 2.82275e-07, 2.821015e-07, 2.823955e-07, 
    2.826766e-07, 2.83148e-07, 2.830704e-07, 2.83278e-07, 2.82388e-07, 
    2.829795e-07, 2.820026e-07, 2.8227e-07, 2.801394e-07, 2.79327e-07, 
    2.789805e-07, 2.786779e-07, 2.779402e-07, 2.784497e-07, 2.782488e-07, 
    2.787267e-07, 2.7903e-07, 2.7888e-07, 2.798053e-07, 2.794457e-07, 
    2.813373e-07, 2.805232e-07, 2.826439e-07, 2.821371e-07, 2.827653e-07, 
    2.824449e-07, 2.829937e-07, 2.824998e-07, 2.833552e-07, 2.835412e-07, 
    2.834141e-07, 2.839026e-07, 2.824724e-07, 2.830219e-07, 2.788758e-07, 
    2.789002e-07, 2.790143e-07, 2.785129e-07, 2.784823e-07, 2.780227e-07, 
    2.784317e-07, 2.786057e-07, 2.790477e-07, 2.793087e-07, 2.795569e-07, 
    2.801021e-07, 2.807103e-07, 2.815601e-07, 2.8217e-07, 2.825784e-07, 
    2.823281e-07, 2.825491e-07, 2.82302e-07, 2.821862e-07, 2.834715e-07, 
    2.8275e-07, 2.838323e-07, 2.837726e-07, 2.832828e-07, 2.837793e-07, 
    2.789174e-07, 2.787767e-07, 2.782874e-07, 2.786703e-07, 2.779726e-07, 
    2.783632e-07, 2.785875e-07, 2.79453e-07, 2.796432e-07, 2.798193e-07, 
    2.801671e-07, 2.80613e-07, 2.813944e-07, 2.820736e-07, 2.82693e-07, 
    2.826477e-07, 2.826636e-07, 2.828019e-07, 2.824593e-07, 2.828581e-07, 
    2.829249e-07, 2.827501e-07, 2.837645e-07, 2.834749e-07, 2.837713e-07, 
    2.835827e-07, 2.788225e-07, 2.790593e-07, 2.789313e-07, 2.791719e-07, 
    2.790024e-07, 2.797558e-07, 2.799815e-07, 2.810368e-07, 2.806041e-07, 
    2.812928e-07, 2.806742e-07, 2.807838e-07, 2.813149e-07, 2.807077e-07, 
    2.820359e-07, 2.811354e-07, 2.828072e-07, 2.819087e-07, 2.828635e-07, 
    2.826904e-07, 2.82977e-07, 2.832336e-07, 2.835563e-07, 2.84151e-07, 
    2.840134e-07, 2.845106e-07, 2.794123e-07, 2.797192e-07, 2.796923e-07, 
    2.800134e-07, 2.802507e-07, 2.80765e-07, 2.815887e-07, 2.812791e-07, 
    2.818475e-07, 2.819614e-07, 2.81098e-07, 2.816281e-07, 2.799246e-07, 
    2.801999e-07, 2.800361e-07, 2.794364e-07, 2.813502e-07, 2.803687e-07, 
    2.8218e-07, 2.816493e-07, 2.83197e-07, 2.824276e-07, 2.839376e-07, 
    2.845814e-07, 2.851875e-07, 2.85894e-07, 2.798868e-07, 2.796783e-07, 
    2.800516e-07, 2.805674e-07, 2.810461e-07, 2.816817e-07, 2.817467e-07, 
    2.818657e-07, 2.821738e-07, 2.824327e-07, 2.819031e-07, 2.824976e-07, 
    2.802634e-07, 2.814354e-07, 2.795993e-07, 2.801525e-07, 2.805371e-07, 
    2.803686e-07, 2.812438e-07, 2.814498e-07, 2.822861e-07, 2.81854e-07, 
    2.844224e-07, 2.832874e-07, 2.86432e-07, 2.855549e-07, 2.796054e-07, 
    2.798861e-07, 2.808617e-07, 2.803978e-07, 2.817241e-07, 2.820501e-07, 
    2.823151e-07, 2.826534e-07, 2.826901e-07, 2.828904e-07, 2.82562e-07, 
    2.828775e-07, 2.81683e-07, 2.822171e-07, 2.807505e-07, 2.811077e-07, 
    2.809435e-07, 2.807631e-07, 2.813195e-07, 2.819114e-07, 2.819243e-07, 
    2.821139e-07, 2.826473e-07, 2.817295e-07, 2.845682e-07, 2.828162e-07, 
    2.80192e-07, 2.807316e-07, 2.80809e-07, 2.806e-07, 2.820174e-07, 
    2.815042e-07, 2.828856e-07, 2.825126e-07, 2.831236e-07, 2.828201e-07, 
    2.827754e-07, 2.823853e-07, 2.821422e-07, 2.815277e-07, 2.810273e-07, 
    2.806304e-07, 2.807227e-07, 2.811587e-07, 2.819476e-07, 2.826932e-07, 
    2.8253e-07, 2.830772e-07, 2.816281e-07, 2.82236e-07, 2.82001e-07, 
    2.826136e-07, 2.812708e-07, 2.824136e-07, 2.809782e-07, 2.811043e-07, 
    2.81494e-07, 2.82277e-07, 2.824505e-07, 2.826353e-07, 2.825213e-07, 
    2.819677e-07, 2.818771e-07, 2.814846e-07, 2.813761e-07, 2.810769e-07, 
    2.808289e-07, 2.810554e-07, 2.812931e-07, 2.819681e-07, 2.825755e-07, 
    2.832371e-07, 2.833991e-07, 2.841703e-07, 2.835422e-07, 2.845779e-07, 
    2.836968e-07, 2.852214e-07, 2.824802e-07, 2.836715e-07, 2.815118e-07, 
    2.817449e-07, 2.82166e-07, 2.831314e-07, 2.826107e-07, 2.832197e-07, 
    2.818735e-07, 2.811736e-07, 2.809927e-07, 2.806544e-07, 2.810004e-07, 
    2.809723e-07, 2.813031e-07, 2.811969e-07, 2.819905e-07, 2.815643e-07, 
    2.827742e-07, 2.83215e-07, 2.844584e-07, 2.852191e-07, 2.859929e-07, 
    2.86334e-07, 2.864378e-07, 2.864812e-07,
  2.756765e-07, 2.764016e-07, 2.762608e-07, 2.768451e-07, 2.765211e-07, 
    2.769035e-07, 2.758237e-07, 2.764303e-07, 2.760432e-07, 2.757419e-07, 
    2.779771e-07, 2.768712e-07, 2.791249e-07, 2.784209e-07, 2.801881e-07, 
    2.790153e-07, 2.804244e-07, 2.801546e-07, 2.80967e-07, 2.807344e-07, 
    2.817716e-07, 2.810743e-07, 2.823091e-07, 2.816053e-07, 2.817154e-07, 
    2.810512e-07, 2.770941e-07, 2.778394e-07, 2.770499e-07, 2.771562e-07, 
    2.771086e-07, 2.765277e-07, 2.762346e-07, 2.756212e-07, 2.757326e-07, 
    2.761833e-07, 2.772041e-07, 2.768579e-07, 2.777304e-07, 2.777107e-07, 
    2.786805e-07, 2.782435e-07, 2.798714e-07, 2.794092e-07, 2.807441e-07, 
    2.804086e-07, 2.807283e-07, 2.806314e-07, 2.807296e-07, 2.802375e-07, 
    2.804483e-07, 2.800153e-07, 2.783253e-07, 2.788224e-07, 2.773386e-07, 
    2.764443e-07, 2.758503e-07, 2.754282e-07, 2.754878e-07, 2.756016e-07, 
    2.761859e-07, 2.767351e-07, 2.771532e-07, 2.774326e-07, 2.777079e-07, 
    2.785398e-07, 2.789802e-07, 2.799647e-07, 2.797874e-07, 2.800879e-07, 
    2.803752e-07, 2.80857e-07, 2.807778e-07, 2.809899e-07, 2.800802e-07, 
    2.806848e-07, 2.796863e-07, 2.799596e-07, 2.777819e-07, 2.769513e-07, 
    2.765973e-07, 2.762878e-07, 2.755337e-07, 2.760545e-07, 2.758493e-07, 
    2.763377e-07, 2.766478e-07, 2.764945e-07, 2.774403e-07, 2.770727e-07, 
    2.790063e-07, 2.781742e-07, 2.803417e-07, 2.798238e-07, 2.804659e-07, 
    2.801384e-07, 2.806993e-07, 2.801945e-07, 2.810689e-07, 2.81259e-07, 
    2.811291e-07, 2.816283e-07, 2.801665e-07, 2.807282e-07, 2.764901e-07, 
    2.765151e-07, 2.766317e-07, 2.761192e-07, 2.760879e-07, 2.756181e-07, 
    2.760362e-07, 2.762141e-07, 2.766658e-07, 2.769327e-07, 2.771863e-07, 
    2.777437e-07, 2.783654e-07, 2.79234e-07, 2.798574e-07, 2.802749e-07, 
    2.80019e-07, 2.802449e-07, 2.799923e-07, 2.798739e-07, 2.811877e-07, 
    2.804503e-07, 2.815566e-07, 2.814954e-07, 2.809949e-07, 2.815023e-07, 
    2.765327e-07, 2.763888e-07, 2.758887e-07, 2.762801e-07, 2.755669e-07, 
    2.759661e-07, 2.761955e-07, 2.770802e-07, 2.772746e-07, 2.774546e-07, 
    2.7781e-07, 2.782658e-07, 2.790646e-07, 2.797588e-07, 2.80392e-07, 
    2.803457e-07, 2.80362e-07, 2.805032e-07, 2.801531e-07, 2.805607e-07, 
    2.80629e-07, 2.804503e-07, 2.814872e-07, 2.811912e-07, 2.814941e-07, 
    2.813014e-07, 2.764356e-07, 2.766777e-07, 2.765469e-07, 2.767929e-07, 
    2.766195e-07, 2.773897e-07, 2.776204e-07, 2.786991e-07, 2.782568e-07, 
    2.789608e-07, 2.783284e-07, 2.784405e-07, 2.789834e-07, 2.783627e-07, 
    2.797204e-07, 2.787999e-07, 2.805087e-07, 2.795904e-07, 2.805662e-07, 
    2.803893e-07, 2.806823e-07, 2.809445e-07, 2.812744e-07, 2.818823e-07, 
    2.817416e-07, 2.822498e-07, 2.770386e-07, 2.773522e-07, 2.773248e-07, 
    2.77653e-07, 2.778956e-07, 2.784212e-07, 2.792632e-07, 2.789467e-07, 
    2.795277e-07, 2.796442e-07, 2.787616e-07, 2.793035e-07, 2.775622e-07, 
    2.778437e-07, 2.776762e-07, 2.770632e-07, 2.790194e-07, 2.780162e-07, 
    2.798676e-07, 2.793251e-07, 2.809071e-07, 2.801207e-07, 2.816641e-07, 
    2.823223e-07, 2.829418e-07, 2.83664e-07, 2.775235e-07, 2.773105e-07, 
    2.77692e-07, 2.782193e-07, 2.787086e-07, 2.793582e-07, 2.794247e-07, 
    2.795463e-07, 2.798613e-07, 2.801259e-07, 2.795846e-07, 2.801922e-07, 
    2.779086e-07, 2.791065e-07, 2.772297e-07, 2.777952e-07, 2.781883e-07, 
    2.780161e-07, 2.789106e-07, 2.791212e-07, 2.799761e-07, 2.795344e-07, 
    2.821598e-07, 2.809996e-07, 2.842139e-07, 2.833173e-07, 2.77236e-07, 
    2.775229e-07, 2.785201e-07, 2.780459e-07, 2.794016e-07, 2.797348e-07, 
    2.800057e-07, 2.803515e-07, 2.803889e-07, 2.805938e-07, 2.802581e-07, 
    2.805806e-07, 2.793596e-07, 2.799055e-07, 2.784064e-07, 2.787716e-07, 
    2.786036e-07, 2.784193e-07, 2.78988e-07, 2.795931e-07, 2.796062e-07, 
    2.798e-07, 2.803454e-07, 2.794071e-07, 2.823088e-07, 2.80518e-07, 
    2.778355e-07, 2.783871e-07, 2.784662e-07, 2.782526e-07, 2.797014e-07, 
    2.791768e-07, 2.805888e-07, 2.802076e-07, 2.808321e-07, 2.805218e-07, 
    2.804762e-07, 2.800774e-07, 2.79829e-07, 2.792008e-07, 2.786894e-07, 
    2.782836e-07, 2.78378e-07, 2.788236e-07, 2.796301e-07, 2.803922e-07, 
    2.802253e-07, 2.807847e-07, 2.793034e-07, 2.799248e-07, 2.796847e-07, 
    2.803108e-07, 2.789383e-07, 2.801064e-07, 2.786392e-07, 2.787681e-07, 
    2.791664e-07, 2.799668e-07, 2.801441e-07, 2.80333e-07, 2.802165e-07, 
    2.796506e-07, 2.79558e-07, 2.791568e-07, 2.790458e-07, 2.7874e-07, 
    2.784866e-07, 2.787181e-07, 2.78961e-07, 2.796509e-07, 2.802719e-07, 
    2.809482e-07, 2.811137e-07, 2.81902e-07, 2.8126e-07, 2.823187e-07, 
    2.814182e-07, 2.829765e-07, 2.801745e-07, 2.813922e-07, 2.791846e-07, 
    2.794229e-07, 2.798534e-07, 2.808401e-07, 2.803079e-07, 2.809304e-07, 
    2.795543e-07, 2.788389e-07, 2.786539e-07, 2.783082e-07, 2.786618e-07, 
    2.786331e-07, 2.789713e-07, 2.788627e-07, 2.796739e-07, 2.792383e-07, 
    2.804749e-07, 2.809255e-07, 2.821965e-07, 2.829741e-07, 2.83765e-07, 
    2.841137e-07, 2.842198e-07, 2.842642e-07,
  2.75814e-07, 2.765496e-07, 2.764067e-07, 2.769995e-07, 2.766708e-07, 
    2.770589e-07, 2.759633e-07, 2.765787e-07, 2.761859e-07, 2.758804e-07, 
    2.781485e-07, 2.77026e-07, 2.793138e-07, 2.785989e-07, 2.803937e-07, 
    2.792025e-07, 2.806337e-07, 2.803596e-07, 2.811849e-07, 2.809485e-07, 
    2.820028e-07, 2.812939e-07, 2.82549e-07, 2.818336e-07, 2.819455e-07, 
    2.812705e-07, 2.772522e-07, 2.780088e-07, 2.772073e-07, 2.773153e-07, 
    2.772669e-07, 2.766775e-07, 2.763802e-07, 2.757579e-07, 2.758709e-07, 
    2.763281e-07, 2.773638e-07, 2.770125e-07, 2.77898e-07, 2.77878e-07, 
    2.788625e-07, 2.784188e-07, 2.800719e-07, 2.796025e-07, 2.809584e-07, 
    2.806176e-07, 2.809423e-07, 2.808439e-07, 2.809436e-07, 2.804437e-07, 
    2.80658e-07, 2.80218e-07, 2.785019e-07, 2.790065e-07, 2.775003e-07, 
    2.765929e-07, 2.759902e-07, 2.755621e-07, 2.756227e-07, 2.75738e-07, 
    2.763308e-07, 2.768878e-07, 2.773121e-07, 2.775957e-07, 2.778751e-07, 
    2.787197e-07, 2.791668e-07, 2.801667e-07, 2.799865e-07, 2.802918e-07, 
    2.805837e-07, 2.810731e-07, 2.809927e-07, 2.812082e-07, 2.802839e-07, 
    2.808982e-07, 2.798838e-07, 2.801614e-07, 2.779504e-07, 2.771073e-07, 
    2.767481e-07, 2.764342e-07, 2.756692e-07, 2.761975e-07, 2.759892e-07, 
    2.764847e-07, 2.767993e-07, 2.766438e-07, 2.776035e-07, 2.772305e-07, 
    2.791933e-07, 2.783484e-07, 2.805496e-07, 2.800235e-07, 2.806757e-07, 
    2.80343e-07, 2.80913e-07, 2.804e-07, 2.812884e-07, 2.814817e-07, 
    2.813496e-07, 2.81857e-07, 2.803716e-07, 2.809423e-07, 2.766394e-07, 
    2.766647e-07, 2.76783e-07, 2.762631e-07, 2.762313e-07, 2.757547e-07, 
    2.761788e-07, 2.763593e-07, 2.768176e-07, 2.770884e-07, 2.773458e-07, 
    2.779114e-07, 2.785426e-07, 2.794245e-07, 2.800576e-07, 2.804817e-07, 
    2.802217e-07, 2.804512e-07, 2.801946e-07, 2.800744e-07, 2.814092e-07, 
    2.806599e-07, 2.817841e-07, 2.817219e-07, 2.812133e-07, 2.817289e-07, 
    2.766826e-07, 2.765366e-07, 2.760292e-07, 2.764263e-07, 2.757028e-07, 
    2.761078e-07, 2.763405e-07, 2.772381e-07, 2.774354e-07, 2.77618e-07, 
    2.779788e-07, 2.784415e-07, 2.792525e-07, 2.799575e-07, 2.806007e-07, 
    2.805536e-07, 2.805702e-07, 2.807137e-07, 2.80358e-07, 2.807721e-07, 
    2.808415e-07, 2.806599e-07, 2.817136e-07, 2.814127e-07, 2.817206e-07, 
    2.815247e-07, 2.76584e-07, 2.768297e-07, 2.766969e-07, 2.769465e-07, 
    2.767706e-07, 2.775522e-07, 2.777864e-07, 2.788814e-07, 2.784323e-07, 
    2.791471e-07, 2.78505e-07, 2.786188e-07, 2.791701e-07, 2.785398e-07, 
    2.799185e-07, 2.789838e-07, 2.807193e-07, 2.797865e-07, 2.807777e-07, 
    2.805979e-07, 2.808956e-07, 2.81162e-07, 2.814973e-07, 2.821152e-07, 
    2.819722e-07, 2.824888e-07, 2.771959e-07, 2.775142e-07, 2.774863e-07, 
    2.778194e-07, 2.780656e-07, 2.785992e-07, 2.794541e-07, 2.791328e-07, 
    2.797227e-07, 2.798411e-07, 2.789448e-07, 2.794951e-07, 2.777273e-07, 
    2.78013e-07, 2.77843e-07, 2.772209e-07, 2.792067e-07, 2.781881e-07, 
    2.80068e-07, 2.795171e-07, 2.81124e-07, 2.803251e-07, 2.818934e-07, 
    2.825625e-07, 2.831923e-07, 2.839269e-07, 2.77688e-07, 2.774717e-07, 
    2.77859e-07, 2.783943e-07, 2.78891e-07, 2.795506e-07, 2.796182e-07, 
    2.797416e-07, 2.800615e-07, 2.803303e-07, 2.797806e-07, 2.803977e-07, 
    2.78079e-07, 2.792951e-07, 2.773899e-07, 2.779638e-07, 2.783628e-07, 
    2.781879e-07, 2.790961e-07, 2.793099e-07, 2.801782e-07, 2.797296e-07, 
    2.823973e-07, 2.812181e-07, 2.844862e-07, 2.835743e-07, 2.773961e-07, 
    2.776873e-07, 2.786996e-07, 2.782182e-07, 2.795947e-07, 2.799331e-07, 
    2.802082e-07, 2.805596e-07, 2.805976e-07, 2.808057e-07, 2.804646e-07, 
    2.807922e-07, 2.79552e-07, 2.801065e-07, 2.785842e-07, 2.789549e-07, 
    2.787844e-07, 2.785973e-07, 2.791747e-07, 2.797892e-07, 2.798025e-07, 
    2.799994e-07, 2.805536e-07, 2.796003e-07, 2.82549e-07, 2.807289e-07, 
    2.780047e-07, 2.785647e-07, 2.786449e-07, 2.78428e-07, 2.798992e-07, 
    2.793664e-07, 2.808006e-07, 2.804133e-07, 2.810479e-07, 2.807326e-07, 
    2.806862e-07, 2.802811e-07, 2.800287e-07, 2.793908e-07, 2.788715e-07, 
    2.784595e-07, 2.785553e-07, 2.790078e-07, 2.798268e-07, 2.806009e-07, 
    2.804314e-07, 2.809997e-07, 2.79495e-07, 2.801262e-07, 2.798822e-07, 
    2.805182e-07, 2.791242e-07, 2.803108e-07, 2.788205e-07, 2.789513e-07, 
    2.793559e-07, 2.801688e-07, 2.803489e-07, 2.805407e-07, 2.804224e-07, 
    2.798476e-07, 2.797535e-07, 2.793461e-07, 2.792334e-07, 2.789229e-07, 
    2.786656e-07, 2.789006e-07, 2.791473e-07, 2.798479e-07, 2.804787e-07, 
    2.811658e-07, 2.81334e-07, 2.821353e-07, 2.814828e-07, 2.825591e-07, 
    2.816437e-07, 2.832278e-07, 2.803798e-07, 2.816171e-07, 2.793743e-07, 
    2.796163e-07, 2.800536e-07, 2.81056e-07, 2.805152e-07, 2.811477e-07, 
    2.797498e-07, 2.790233e-07, 2.788355e-07, 2.784845e-07, 2.788435e-07, 
    2.788143e-07, 2.791577e-07, 2.790474e-07, 2.798712e-07, 2.794288e-07, 
    2.80685e-07, 2.811428e-07, 2.824346e-07, 2.832252e-07, 2.840296e-07, 
    2.843843e-07, 2.844922e-07, 2.845374e-07,
  2.694084e-07, 2.701424e-07, 2.699998e-07, 2.705915e-07, 2.702633e-07, 
    2.706507e-07, 2.695573e-07, 2.701715e-07, 2.697794e-07, 2.694746e-07, 
    2.717391e-07, 2.706179e-07, 2.729035e-07, 2.72189e-07, 2.739836e-07, 
    2.727923e-07, 2.742237e-07, 2.739494e-07, 2.747753e-07, 2.745387e-07, 
    2.755944e-07, 2.748845e-07, 2.761416e-07, 2.75425e-07, 2.75537e-07, 
    2.74861e-07, 2.708437e-07, 2.715996e-07, 2.707989e-07, 2.709067e-07, 
    2.708584e-07, 2.7027e-07, 2.699734e-07, 2.693524e-07, 2.694651e-07, 
    2.699213e-07, 2.709552e-07, 2.706044e-07, 2.714886e-07, 2.714687e-07, 
    2.724524e-07, 2.720089e-07, 2.736616e-07, 2.731921e-07, 2.745486e-07, 
    2.742076e-07, 2.745326e-07, 2.744341e-07, 2.745338e-07, 2.740337e-07, 
    2.74248e-07, 2.738078e-07, 2.72092e-07, 2.725964e-07, 2.710915e-07, 
    2.701858e-07, 2.695842e-07, 2.691571e-07, 2.692175e-07, 2.693326e-07, 
    2.69924e-07, 2.704799e-07, 2.709035e-07, 2.711867e-07, 2.714658e-07, 
    2.723098e-07, 2.727567e-07, 2.737565e-07, 2.735762e-07, 2.738817e-07, 
    2.741736e-07, 2.746635e-07, 2.745829e-07, 2.747987e-07, 2.738737e-07, 
    2.744885e-07, 2.734735e-07, 2.737511e-07, 2.715412e-07, 2.706991e-07, 
    2.703406e-07, 2.700272e-07, 2.692639e-07, 2.69791e-07, 2.695832e-07, 
    2.700775e-07, 2.703916e-07, 2.702363e-07, 2.711945e-07, 2.70822e-07, 
    2.727831e-07, 2.719387e-07, 2.741396e-07, 2.736132e-07, 2.742657e-07, 
    2.739328e-07, 2.745032e-07, 2.739899e-07, 2.74879e-07, 2.750725e-07, 
    2.749403e-07, 2.754483e-07, 2.739614e-07, 2.745325e-07, 2.702319e-07, 
    2.702572e-07, 2.703752e-07, 2.698564e-07, 2.698247e-07, 2.693492e-07, 
    2.697724e-07, 2.699525e-07, 2.704098e-07, 2.706801e-07, 2.709371e-07, 
    2.71502e-07, 2.721327e-07, 2.730142e-07, 2.736473e-07, 2.740715e-07, 
    2.738115e-07, 2.740411e-07, 2.737844e-07, 2.736641e-07, 2.75e-07, 
    2.742499e-07, 2.753752e-07, 2.75313e-07, 2.748038e-07, 2.7532e-07, 
    2.70275e-07, 2.701293e-07, 2.696231e-07, 2.700193e-07, 2.692975e-07, 
    2.697015e-07, 2.699337e-07, 2.708297e-07, 2.710266e-07, 2.71209e-07, 
    2.715693e-07, 2.720316e-07, 2.728422e-07, 2.735472e-07, 2.741906e-07, 
    2.741435e-07, 2.741601e-07, 2.743037e-07, 2.739478e-07, 2.743622e-07, 
    2.744317e-07, 2.742499e-07, 2.753047e-07, 2.750034e-07, 2.753117e-07, 
    2.751156e-07, 2.701767e-07, 2.704219e-07, 2.702894e-07, 2.705385e-07, 
    2.70363e-07, 2.711433e-07, 2.713772e-07, 2.724713e-07, 2.720225e-07, 
    2.727369e-07, 2.720951e-07, 2.722088e-07, 2.7276e-07, 2.721298e-07, 
    2.735083e-07, 2.725737e-07, 2.743093e-07, 2.733764e-07, 2.743677e-07, 
    2.741878e-07, 2.744858e-07, 2.747525e-07, 2.750881e-07, 2.75707e-07, 
    2.755637e-07, 2.760812e-07, 2.707874e-07, 2.711053e-07, 2.710774e-07, 
    2.714101e-07, 2.716561e-07, 2.721892e-07, 2.730438e-07, 2.727225e-07, 
    2.733124e-07, 2.734307e-07, 2.725346e-07, 2.730848e-07, 2.713181e-07, 
    2.716036e-07, 2.714337e-07, 2.708125e-07, 2.727964e-07, 2.717785e-07, 
    2.736578e-07, 2.731067e-07, 2.747144e-07, 2.73915e-07, 2.754848e-07, 
    2.761552e-07, 2.767862e-07, 2.77523e-07, 2.712789e-07, 2.710629e-07, 
    2.714497e-07, 2.719845e-07, 2.724809e-07, 2.731403e-07, 2.732078e-07, 
    2.733313e-07, 2.736512e-07, 2.739201e-07, 2.733703e-07, 2.739875e-07, 
    2.716697e-07, 2.728848e-07, 2.709812e-07, 2.715545e-07, 2.71953e-07, 
    2.717783e-07, 2.726858e-07, 2.728996e-07, 2.73768e-07, 2.733192e-07, 
    2.759897e-07, 2.748087e-07, 2.780839e-07, 2.771693e-07, 2.709874e-07, 
    2.712782e-07, 2.722896e-07, 2.718085e-07, 2.731844e-07, 2.735228e-07, 
    2.73798e-07, 2.741495e-07, 2.741875e-07, 2.743958e-07, 2.740545e-07, 
    2.743823e-07, 2.731417e-07, 2.736963e-07, 2.721742e-07, 2.725447e-07, 
    2.723743e-07, 2.721873e-07, 2.727644e-07, 2.733789e-07, 2.733922e-07, 
    2.735891e-07, 2.741438e-07, 2.7319e-07, 2.761418e-07, 2.743193e-07, 
    2.715952e-07, 2.721548e-07, 2.722349e-07, 2.720181e-07, 2.734889e-07, 
    2.729561e-07, 2.743907e-07, 2.740032e-07, 2.746382e-07, 2.743226e-07, 
    2.742762e-07, 2.738709e-07, 2.736184e-07, 2.729805e-07, 2.724613e-07, 
    2.720496e-07, 2.721453e-07, 2.725976e-07, 2.734165e-07, 2.741909e-07, 
    2.740213e-07, 2.745899e-07, 2.730847e-07, 2.73716e-07, 2.73472e-07, 
    2.741081e-07, 2.727139e-07, 2.739009e-07, 2.724104e-07, 2.725411e-07, 
    2.729456e-07, 2.737587e-07, 2.739387e-07, 2.741307e-07, 2.740122e-07, 
    2.734373e-07, 2.733432e-07, 2.729358e-07, 2.728232e-07, 2.725127e-07, 
    2.722555e-07, 2.724904e-07, 2.727371e-07, 2.734376e-07, 2.740686e-07, 
    2.747562e-07, 2.749246e-07, 2.757273e-07, 2.750737e-07, 2.761519e-07, 
    2.752351e-07, 2.76822e-07, 2.739698e-07, 2.752083e-07, 2.72964e-07, 
    2.73206e-07, 2.736434e-07, 2.746465e-07, 2.741051e-07, 2.747382e-07, 
    2.733395e-07, 2.726132e-07, 2.724253e-07, 2.720746e-07, 2.724333e-07, 
    2.724042e-07, 2.727474e-07, 2.726371e-07, 2.734609e-07, 2.730185e-07, 
    2.74275e-07, 2.747333e-07, 2.760269e-07, 2.768193e-07, 2.776258e-07, 
    2.779816e-07, 2.780899e-07, 2.781352e-07,
  2.510149e-07, 2.517251e-07, 2.51587e-07, 2.521599e-07, 2.518421e-07, 
    2.522173e-07, 2.511589e-07, 2.517532e-07, 2.513738e-07, 2.510789e-07, 
    2.532723e-07, 2.521855e-07, 2.54402e-07, 2.537084e-07, 2.554515e-07, 
    2.542941e-07, 2.55685e-07, 2.554182e-07, 2.562215e-07, 2.559914e-07, 
    2.570194e-07, 2.563278e-07, 2.575525e-07, 2.568542e-07, 2.569634e-07, 
    2.56305e-07, 2.524042e-07, 2.53137e-07, 2.523608e-07, 2.524652e-07, 
    2.524183e-07, 2.518487e-07, 2.515616e-07, 2.509607e-07, 2.510698e-07, 
    2.515112e-07, 2.525122e-07, 2.521724e-07, 2.530291e-07, 2.530097e-07, 
    2.53964e-07, 2.535337e-07, 2.551384e-07, 2.546822e-07, 2.56001e-07, 
    2.556692e-07, 2.559854e-07, 2.558895e-07, 2.559866e-07, 2.555001e-07, 
    2.557085e-07, 2.552805e-07, 2.536142e-07, 2.541038e-07, 2.526442e-07, 
    2.517672e-07, 2.511849e-07, 2.507719e-07, 2.508303e-07, 2.509416e-07, 
    2.515137e-07, 2.520518e-07, 2.524621e-07, 2.527365e-07, 2.53007e-07, 
    2.538258e-07, 2.542594e-07, 2.552307e-07, 2.550554e-07, 2.553524e-07, 
    2.556362e-07, 2.561128e-07, 2.560343e-07, 2.562443e-07, 2.553446e-07, 
    2.559425e-07, 2.549555e-07, 2.552254e-07, 2.530804e-07, 2.52264e-07, 
    2.519171e-07, 2.516135e-07, 2.508752e-07, 2.51385e-07, 2.51184e-07, 
    2.516623e-07, 2.519662e-07, 2.518159e-07, 2.52744e-07, 2.523831e-07, 
    2.542851e-07, 2.534656e-07, 2.556031e-07, 2.550914e-07, 2.557258e-07, 
    2.55402e-07, 2.559568e-07, 2.554575e-07, 2.563225e-07, 2.565109e-07, 
    2.563822e-07, 2.568769e-07, 2.554298e-07, 2.559854e-07, 2.518117e-07, 
    2.518362e-07, 2.519504e-07, 2.514484e-07, 2.514176e-07, 2.509577e-07, 
    2.51367e-07, 2.515413e-07, 2.519839e-07, 2.522457e-07, 2.524947e-07, 
    2.530421e-07, 2.536538e-07, 2.545095e-07, 2.551245e-07, 2.555369e-07, 
    2.55284e-07, 2.555073e-07, 2.552577e-07, 2.551407e-07, 2.564403e-07, 
    2.557105e-07, 2.568057e-07, 2.567451e-07, 2.562493e-07, 2.567519e-07, 
    2.518534e-07, 2.517124e-07, 2.512226e-07, 2.516059e-07, 2.509076e-07, 
    2.512984e-07, 2.515231e-07, 2.523906e-07, 2.525813e-07, 2.527581e-07, 
    2.531074e-07, 2.535557e-07, 2.543424e-07, 2.550273e-07, 2.556527e-07, 
    2.556069e-07, 2.55623e-07, 2.557628e-07, 2.554166e-07, 2.558196e-07, 
    2.558872e-07, 2.557104e-07, 2.567369e-07, 2.564436e-07, 2.567438e-07, 
    2.565528e-07, 2.517582e-07, 2.519956e-07, 2.518673e-07, 2.521086e-07, 
    2.519386e-07, 2.526945e-07, 2.529212e-07, 2.539824e-07, 2.535469e-07, 
    2.542402e-07, 2.536173e-07, 2.537276e-07, 2.542628e-07, 2.536509e-07, 
    2.549895e-07, 2.540819e-07, 2.557682e-07, 2.548614e-07, 2.55825e-07, 
    2.5565e-07, 2.559398e-07, 2.561994e-07, 2.565261e-07, 2.571289e-07, 
    2.569893e-07, 2.574936e-07, 2.523496e-07, 2.526577e-07, 2.526306e-07, 
    2.52953e-07, 2.531915e-07, 2.537085e-07, 2.545382e-07, 2.542262e-07, 
    2.54799e-07, 2.54914e-07, 2.540438e-07, 2.54578e-07, 2.528639e-07, 
    2.531407e-07, 2.529759e-07, 2.523739e-07, 2.54298e-07, 2.533103e-07, 
    2.551347e-07, 2.545993e-07, 2.561624e-07, 2.553848e-07, 2.569124e-07, 
    2.575659e-07, 2.581812e-07, 2.589006e-07, 2.528258e-07, 2.526165e-07, 
    2.529914e-07, 2.535101e-07, 2.539916e-07, 2.546319e-07, 2.546975e-07, 
    2.548174e-07, 2.551283e-07, 2.553897e-07, 2.548554e-07, 2.554552e-07, 
    2.532049e-07, 2.543838e-07, 2.525373e-07, 2.530931e-07, 2.534795e-07, 
    2.5331e-07, 2.541905e-07, 2.543981e-07, 2.552419e-07, 2.548056e-07, 
    2.574046e-07, 2.562542e-07, 2.594486e-07, 2.585552e-07, 2.525434e-07, 
    2.528251e-07, 2.538061e-07, 2.533393e-07, 2.546747e-07, 2.550035e-07, 
    2.552709e-07, 2.556128e-07, 2.556497e-07, 2.558523e-07, 2.555203e-07, 
    2.558392e-07, 2.546333e-07, 2.551721e-07, 2.536939e-07, 2.540536e-07, 
    2.538881e-07, 2.537067e-07, 2.542668e-07, 2.548637e-07, 2.548765e-07, 
    2.55068e-07, 2.556076e-07, 2.546801e-07, 2.575531e-07, 2.557782e-07, 
    2.531324e-07, 2.536753e-07, 2.537529e-07, 2.535426e-07, 2.549706e-07, 
    2.54453e-07, 2.558474e-07, 2.554704e-07, 2.560881e-07, 2.557811e-07, 
    2.55736e-07, 2.553418e-07, 2.550964e-07, 2.544767e-07, 2.539727e-07, 
    2.535731e-07, 2.53666e-07, 2.541049e-07, 2.549003e-07, 2.55653e-07, 
    2.554881e-07, 2.560411e-07, 2.545778e-07, 2.551913e-07, 2.549541e-07, 
    2.555725e-07, 2.542179e-07, 2.553713e-07, 2.539232e-07, 2.540501e-07, 
    2.544427e-07, 2.552328e-07, 2.554077e-07, 2.555944e-07, 2.554792e-07, 
    2.549205e-07, 2.54829e-07, 2.544332e-07, 2.543239e-07, 2.540224e-07, 
    2.537729e-07, 2.540009e-07, 2.542404e-07, 2.549207e-07, 2.555341e-07, 
    2.562031e-07, 2.563669e-07, 2.571489e-07, 2.565122e-07, 2.57563e-07, 
    2.566696e-07, 2.582165e-07, 2.554382e-07, 2.566433e-07, 2.544606e-07, 
    2.546956e-07, 2.551208e-07, 2.560963e-07, 2.555696e-07, 2.561856e-07, 
    2.548254e-07, 2.541201e-07, 2.539377e-07, 2.535974e-07, 2.539455e-07, 
    2.539172e-07, 2.542503e-07, 2.541432e-07, 2.549433e-07, 2.545135e-07, 
    2.557348e-07, 2.561808e-07, 2.574407e-07, 2.582136e-07, 2.590009e-07, 
    2.593486e-07, 2.594544e-07, 2.594986e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  7.623649e-08, 7.644516e-08, 7.640461e-08, 7.657286e-08, 7.647954e-08, 
    7.658971e-08, 7.627882e-08, 7.645342e-08, 7.634197e-08, 7.62553e-08, 
    7.689925e-08, 7.658038e-08, 7.723048e-08, 7.70272e-08, 7.753781e-08, 
    7.719884e-08, 7.760615e-08, 7.752807e-08, 7.776314e-08, 7.76958e-08, 
    7.799632e-08, 7.779421e-08, 7.815211e-08, 7.794808e-08, 7.797998e-08, 
    7.778754e-08, 7.664459e-08, 7.685954e-08, 7.663184e-08, 7.66625e-08, 
    7.664875e-08, 7.648146e-08, 7.639712e-08, 7.622056e-08, 7.625263e-08, 
    7.638231e-08, 7.667629e-08, 7.657653e-08, 7.682798e-08, 7.682231e-08, 
    7.710213e-08, 7.697598e-08, 7.744618e-08, 7.731258e-08, 7.769862e-08, 
    7.760154e-08, 7.769405e-08, 7.766601e-08, 7.769442e-08, 7.755205e-08, 
    7.761304e-08, 7.748777e-08, 7.69996e-08, 7.714308e-08, 7.671504e-08, 
    7.64575e-08, 7.628647e-08, 7.616506e-08, 7.618222e-08, 7.621494e-08, 
    7.638307e-08, 7.654115e-08, 7.666159e-08, 7.674213e-08, 7.682149e-08, 
    7.706157e-08, 7.718869e-08, 7.747317e-08, 7.742187e-08, 7.750881e-08, 
    7.759189e-08, 7.773131e-08, 7.770838e-08, 7.776979e-08, 7.750653e-08, 
    7.768149e-08, 7.739264e-08, 7.747165e-08, 7.684295e-08, 7.660345e-08, 
    7.650154e-08, 7.64124e-08, 7.619542e-08, 7.634526e-08, 7.628619e-08, 
    7.642673e-08, 7.651601e-08, 7.647186e-08, 7.674434e-08, 7.663841e-08, 
    7.719622e-08, 7.695601e-08, 7.758219e-08, 7.74324e-08, 7.76181e-08, 
    7.752336e-08, 7.768568e-08, 7.75396e-08, 7.779266e-08, 7.784774e-08, 
    7.781009e-08, 7.795472e-08, 7.753149e-08, 7.769404e-08, 7.647062e-08, 
    7.647782e-08, 7.651137e-08, 7.636387e-08, 7.635484e-08, 7.621968e-08, 
    7.633997e-08, 7.639117e-08, 7.65212e-08, 7.659807e-08, 7.667116e-08, 
    7.683181e-08, 7.701119e-08, 7.726197e-08, 7.744212e-08, 7.756284e-08, 
    7.748882e-08, 7.755416e-08, 7.748111e-08, 7.744688e-08, 7.782709e-08, 
    7.761361e-08, 7.793392e-08, 7.791621e-08, 7.777125e-08, 7.791819e-08, 
    7.648288e-08, 7.644144e-08, 7.629752e-08, 7.641015e-08, 7.620496e-08, 
    7.631981e-08, 7.638584e-08, 7.66406e-08, 7.669659e-08, 7.674847e-08, 
    7.685095e-08, 7.698243e-08, 7.721304e-08, 7.741363e-08, 7.759672e-08, 
    7.758331e-08, 7.758803e-08, 7.762892e-08, 7.752763e-08, 7.764555e-08, 
    7.766533e-08, 7.76136e-08, 7.791383e-08, 7.782807e-08, 7.791583e-08, 
    7.785999e-08, 7.645492e-08, 7.652464e-08, 7.648696e-08, 7.65578e-08, 
    7.650789e-08, 7.672979e-08, 7.679631e-08, 7.710752e-08, 7.697984e-08, 
    7.718307e-08, 7.700049e-08, 7.703284e-08, 7.718965e-08, 7.701037e-08, 
    7.740255e-08, 7.713665e-08, 7.76305e-08, 7.736501e-08, 7.764714e-08, 
    7.759594e-08, 7.768072e-08, 7.775665e-08, 7.785217e-08, 7.802836e-08, 
    7.798757e-08, 7.813491e-08, 7.662858e-08, 7.671898e-08, 7.671105e-08, 
    7.680566e-08, 7.687562e-08, 7.702726e-08, 7.727039e-08, 7.717897e-08, 
    7.73468e-08, 7.738048e-08, 7.712552e-08, 7.728205e-08, 7.67795e-08, 
    7.686069e-08, 7.681236e-08, 7.66357e-08, 7.720001e-08, 7.691045e-08, 
    7.744509e-08, 7.728828e-08, 7.774582e-08, 7.751829e-08, 7.796511e-08, 
    7.815598e-08, 7.833569e-08, 7.854553e-08, 7.676834e-08, 7.670692e-08, 
    7.681692e-08, 7.696904e-08, 7.711023e-08, 7.729785e-08, 7.731705e-08, 
    7.735219e-08, 7.744323e-08, 7.751974e-08, 7.736328e-08, 7.753892e-08, 
    7.687949e-08, 7.722515e-08, 7.668368e-08, 7.684673e-08, 7.696008e-08, 
    7.691038e-08, 7.716854e-08, 7.722935e-08, 7.747646e-08, 7.734874e-08, 
    7.810886e-08, 7.777265e-08, 7.870533e-08, 7.844478e-08, 7.668545e-08, 
    7.676814e-08, 7.705584e-08, 7.691897e-08, 7.731038e-08, 7.740669e-08, 
    7.748498e-08, 7.758503e-08, 7.759585e-08, 7.765512e-08, 7.755798e-08, 
    7.765129e-08, 7.729825e-08, 7.745604e-08, 7.702298e-08, 7.71284e-08, 
    7.707991e-08, 7.702671e-08, 7.71909e-08, 7.736573e-08, 7.736951e-08, 
    7.742555e-08, 7.758342e-08, 7.731197e-08, 7.815218e-08, 7.763335e-08, 
    7.68583e-08, 7.701748e-08, 7.704026e-08, 7.697859e-08, 7.739703e-08, 
    7.724544e-08, 7.765367e-08, 7.754338e-08, 7.77241e-08, 7.76343e-08, 
    7.762108e-08, 7.750573e-08, 7.74339e-08, 7.725239e-08, 7.710467e-08, 
    7.698755e-08, 7.701478e-08, 7.714345e-08, 7.737644e-08, 7.759681e-08, 
    7.754854e-08, 7.771037e-08, 7.728201e-08, 7.746164e-08, 7.739221e-08, 
    7.757325e-08, 7.717654e-08, 7.751427e-08, 7.709018e-08, 7.712737e-08, 
    7.724243e-08, 7.74738e-08, 7.752503e-08, 7.757966e-08, 7.754596e-08, 
    7.738236e-08, 7.735557e-08, 7.723964e-08, 7.720762e-08, 7.711928e-08, 
    7.704612e-08, 7.711296e-08, 7.718313e-08, 7.738244e-08, 7.7562e-08, 
    7.775772e-08, 7.780563e-08, 7.803415e-08, 7.784809e-08, 7.815506e-08, 
    7.789401e-08, 7.834588e-08, 7.753389e-08, 7.788639e-08, 7.724768e-08, 
    7.731652e-08, 7.744099e-08, 7.772646e-08, 7.757239e-08, 7.775259e-08, 
    7.735452e-08, 7.714787e-08, 7.709443e-08, 7.699466e-08, 7.709671e-08, 
    7.708842e-08, 7.718606e-08, 7.715469e-08, 7.738906e-08, 7.726317e-08, 
    7.762075e-08, 7.775118e-08, 7.811946e-08, 7.834512e-08, 7.857481e-08, 
    7.867618e-08, 7.870703e-08, 7.871993e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.949716e-13, 9.975021e-13, 9.970106e-13, 9.990496e-13, 9.979191e-13, 
    9.992536e-13, 9.954853e-13, 9.976022e-13, 9.962513e-13, 9.952001e-13, 
    1.003e-12, 9.991407e-13, 1.007005e-12, 1.004549e-12, 1.010716e-12, 
    1.006623e-12, 1.01154e-12, 1.010599e-12, 1.013433e-12, 1.012622e-12, 
    1.016241e-12, 1.013808e-12, 1.018117e-12, 1.015661e-12, 1.016045e-12, 
    1.013728e-12, 9.999188e-13, 1.00252e-12, 9.997643e-13, 1.000136e-12, 
    9.999692e-13, 9.979422e-13, 9.969193e-13, 9.947787e-13, 9.951677e-13, 
    9.967402e-13, 1.000302e-12, 9.990944e-13, 1.002139e-12, 1.002071e-12, 
    1.005455e-12, 1.00393e-12, 1.009611e-12, 1.007998e-12, 1.012656e-12, 
    1.011485e-12, 1.012601e-12, 1.012263e-12, 1.012605e-12, 1.010888e-12, 
    1.011624e-12, 1.010113e-12, 1.004215e-12, 1.00595e-12, 1.000772e-12, 
    9.97651e-13, 9.955781e-13, 9.941052e-13, 9.943135e-13, 9.947103e-13, 
    9.967493e-13, 9.986657e-13, 1.000125e-12, 1.0011e-12, 1.002061e-12, 
    1.004964e-12, 1.0065e-12, 1.009936e-12, 1.009317e-12, 1.010366e-12, 
    1.011369e-12, 1.01305e-12, 1.012773e-12, 1.013513e-12, 1.010339e-12, 
    1.012449e-12, 1.008965e-12, 1.009918e-12, 1.002319e-12, 9.994205e-13, 
    9.981848e-13, 9.971051e-13, 9.944735e-13, 9.962909e-13, 9.955746e-13, 
    9.972791e-13, 9.983611e-13, 9.978262e-13, 1.001127e-12, 9.99844e-13, 
    1.006592e-12, 1.003688e-12, 1.011252e-12, 1.009444e-12, 1.011685e-12, 
    1.010542e-12, 1.0125e-12, 1.010738e-12, 1.013789e-12, 1.014453e-12, 
    1.013999e-12, 1.015741e-12, 1.01064e-12, 1.0126e-12, 9.97811e-13, 
    9.978983e-13, 9.98305e-13, 9.965165e-13, 9.964073e-13, 9.947679e-13, 
    9.96227e-13, 9.968477e-13, 9.98424e-13, 9.993553e-13, 1.00024e-12, 
    1.002185e-12, 1.004355e-12, 1.007386e-12, 1.009562e-12, 1.011018e-12, 
    1.010125e-12, 1.010914e-12, 1.010032e-12, 1.009619e-12, 1.014204e-12, 
    1.01163e-12, 1.015491e-12, 1.015278e-12, 1.013531e-12, 1.015302e-12, 
    9.979595e-13, 9.974574e-13, 9.957122e-13, 9.970781e-13, 9.945893e-13, 
    9.959824e-13, 9.967827e-13, 9.998701e-13, 1.000549e-12, 1.001177e-12, 
    1.002417e-12, 1.004008e-12, 1.006795e-12, 1.009218e-12, 1.011427e-12, 
    1.011265e-12, 1.011322e-12, 1.011815e-12, 1.010594e-12, 1.012016e-12, 
    1.012254e-12, 1.011631e-12, 1.015249e-12, 1.014216e-12, 1.015273e-12, 
    1.014601e-12, 9.976207e-13, 9.984656e-13, 9.980091e-13, 9.988674e-13, 
    9.982625e-13, 1.00095e-12, 1.001755e-12, 1.00552e-12, 1.003976e-12, 
    1.006433e-12, 1.004226e-12, 1.004617e-12, 1.006512e-12, 1.004346e-12, 
    1.009083e-12, 1.005871e-12, 1.011834e-12, 1.00863e-12, 1.012035e-12, 
    1.011418e-12, 1.01244e-12, 1.013355e-12, 1.014506e-12, 1.016628e-12, 
    1.016137e-12, 1.01791e-12, 9.997249e-13, 1.000819e-12, 1.000724e-12, 
    1.001869e-12, 1.002715e-12, 1.00455e-12, 1.007488e-12, 1.006384e-12, 
    1.008411e-12, 1.008818e-12, 1.005738e-12, 1.007629e-12, 1.001552e-12, 
    1.002534e-12, 1.00195e-12, 9.99811e-13, 1.006637e-12, 1.003136e-12, 
    1.009597e-12, 1.007704e-12, 1.013225e-12, 1.01048e-12, 1.015866e-12, 
    1.018163e-12, 1.020324e-12, 1.022845e-12, 1.001417e-12, 1.000674e-12, 
    1.002005e-12, 1.003845e-12, 1.005553e-12, 1.00782e-12, 1.008052e-12, 
    1.008476e-12, 1.009575e-12, 1.010498e-12, 1.00861e-12, 1.01073e-12, 
    1.002761e-12, 1.006941e-12, 1.000392e-12, 1.002366e-12, 1.003737e-12, 
    1.003136e-12, 1.006258e-12, 1.006993e-12, 1.009976e-12, 1.008434e-12, 
    1.017596e-12, 1.013548e-12, 1.024763e-12, 1.021635e-12, 1.000414e-12, 
    1.001415e-12, 1.004895e-12, 1.00324e-12, 1.007971e-12, 1.009134e-12, 
    1.010079e-12, 1.011286e-12, 1.011416e-12, 1.012131e-12, 1.01096e-12, 
    1.012085e-12, 1.007824e-12, 1.00973e-12, 1.004498e-12, 1.005772e-12, 
    1.005186e-12, 1.004543e-12, 1.006528e-12, 1.008639e-12, 1.008685e-12, 
    1.009362e-12, 1.011265e-12, 1.00799e-12, 1.018116e-12, 1.011867e-12, 
    1.002506e-12, 1.004431e-12, 1.004707e-12, 1.003961e-12, 1.009017e-12, 
    1.007187e-12, 1.012114e-12, 1.010784e-12, 1.012963e-12, 1.01188e-12, 
    1.011721e-12, 1.010329e-12, 1.009462e-12, 1.00727e-12, 1.005486e-12, 
    1.00407e-12, 1.004399e-12, 1.005954e-12, 1.008768e-12, 1.011428e-12, 
    1.010845e-12, 1.012797e-12, 1.007628e-12, 1.009797e-12, 1.008959e-12, 
    1.011144e-12, 1.006354e-12, 1.010431e-12, 1.005311e-12, 1.00576e-12, 
    1.00715e-12, 1.009943e-12, 1.010562e-12, 1.011221e-12, 1.010815e-12, 
    1.00884e-12, 1.008517e-12, 1.007117e-12, 1.00673e-12, 1.005662e-12, 
    1.004778e-12, 1.005586e-12, 1.006434e-12, 1.008841e-12, 1.011008e-12, 
    1.013368e-12, 1.013946e-12, 1.016696e-12, 1.014456e-12, 1.01815e-12, 
    1.015008e-12, 1.020446e-12, 1.010668e-12, 1.014917e-12, 1.007214e-12, 
    1.008045e-12, 1.009548e-12, 1.012991e-12, 1.011134e-12, 1.013306e-12, 
    1.008504e-12, 1.006007e-12, 1.005362e-12, 1.004156e-12, 1.00539e-12, 
    1.005289e-12, 1.006469e-12, 1.00609e-12, 1.008921e-12, 1.007401e-12, 
    1.011717e-12, 1.013289e-12, 1.017724e-12, 1.020437e-12, 1.023197e-12, 
    1.024414e-12, 1.024784e-12, 1.024938e-12 ;

 LITR1C =
  3.066706e-05, 3.066695e-05, 3.066697e-05, 3.066688e-05, 3.066693e-05, 
    3.066687e-05, 3.066704e-05, 3.066694e-05, 3.0667e-05, 3.066705e-05, 
    3.06667e-05, 3.066687e-05, 3.066651e-05, 3.066663e-05, 3.066635e-05, 
    3.066653e-05, 3.066631e-05, 3.066635e-05, 3.066622e-05, 3.066626e-05, 
    3.066609e-05, 3.066621e-05, 3.066601e-05, 3.066612e-05, 3.066611e-05, 
    3.066621e-05, 3.066684e-05, 3.066672e-05, 3.066684e-05, 3.066683e-05, 
    3.066683e-05, 3.066692e-05, 3.066697e-05, 3.066707e-05, 3.066705e-05, 
    3.066698e-05, 3.066682e-05, 3.066687e-05, 3.066674e-05, 3.066674e-05, 
    3.066659e-05, 3.066666e-05, 3.06664e-05, 3.066647e-05, 3.066626e-05, 
    3.066631e-05, 3.066626e-05, 3.066628e-05, 3.066626e-05, 3.066634e-05, 
    3.066631e-05, 3.066638e-05, 3.066664e-05, 3.066656e-05, 3.06668e-05, 
    3.066694e-05, 3.066703e-05, 3.06671e-05, 3.066709e-05, 3.066707e-05, 
    3.066698e-05, 3.066689e-05, 3.066683e-05, 3.066678e-05, 3.066674e-05, 
    3.066661e-05, 3.066654e-05, 3.066638e-05, 3.066641e-05, 3.066636e-05, 
    3.066632e-05, 3.066624e-05, 3.066626e-05, 3.066622e-05, 3.066636e-05, 
    3.066627e-05, 3.066643e-05, 3.066638e-05, 3.066673e-05, 3.066686e-05, 
    3.066691e-05, 3.066696e-05, 3.066708e-05, 3.0667e-05, 3.066703e-05, 
    3.066696e-05, 3.066691e-05, 3.066693e-05, 3.066678e-05, 3.066684e-05, 
    3.066654e-05, 3.066667e-05, 3.066632e-05, 3.06664e-05, 3.06663e-05, 
    3.066635e-05, 3.066627e-05, 3.066635e-05, 3.066621e-05, 3.066618e-05, 
    3.06662e-05, 3.066612e-05, 3.066635e-05, 3.066626e-05, 3.066693e-05, 
    3.066693e-05, 3.066691e-05, 3.066699e-05, 3.066699e-05, 3.066707e-05, 
    3.0667e-05, 3.066698e-05, 3.06669e-05, 3.066686e-05, 3.066682e-05, 
    3.066673e-05, 3.066663e-05, 3.06665e-05, 3.06664e-05, 3.066633e-05, 
    3.066638e-05, 3.066634e-05, 3.066638e-05, 3.06664e-05, 3.066619e-05, 
    3.066631e-05, 3.066613e-05, 3.066614e-05, 3.066622e-05, 3.066614e-05, 
    3.066692e-05, 3.066695e-05, 3.066703e-05, 3.066696e-05, 3.066708e-05, 
    3.066702e-05, 3.066698e-05, 3.066684e-05, 3.066681e-05, 3.066678e-05, 
    3.066672e-05, 3.066665e-05, 3.066652e-05, 3.066642e-05, 3.066631e-05, 
    3.066632e-05, 3.066632e-05, 3.06663e-05, 3.066635e-05, 3.066629e-05, 
    3.066628e-05, 3.066631e-05, 3.066614e-05, 3.066619e-05, 3.066614e-05, 
    3.066617e-05, 3.066694e-05, 3.06669e-05, 3.066692e-05, 3.066688e-05, 
    3.066691e-05, 3.066679e-05, 3.066675e-05, 3.066658e-05, 3.066665e-05, 
    3.066654e-05, 3.066664e-05, 3.066662e-05, 3.066654e-05, 3.066664e-05, 
    3.066642e-05, 3.066657e-05, 3.06663e-05, 3.066644e-05, 3.066629e-05, 
    3.066632e-05, 3.066627e-05, 3.066623e-05, 3.066618e-05, 3.066608e-05, 
    3.06661e-05, 3.066602e-05, 3.066684e-05, 3.06668e-05, 3.06668e-05, 
    3.066675e-05, 3.066671e-05, 3.066663e-05, 3.066649e-05, 3.066654e-05, 
    3.066645e-05, 3.066643e-05, 3.066657e-05, 3.066649e-05, 3.066676e-05, 
    3.066672e-05, 3.066674e-05, 3.066684e-05, 3.066653e-05, 3.066669e-05, 
    3.06664e-05, 3.066648e-05, 3.066623e-05, 3.066636e-05, 3.066611e-05, 
    3.066601e-05, 3.066591e-05, 3.06658e-05, 3.066677e-05, 3.06668e-05, 
    3.066674e-05, 3.066666e-05, 3.066658e-05, 3.066648e-05, 3.066647e-05, 
    3.066645e-05, 3.06664e-05, 3.066636e-05, 3.066644e-05, 3.066635e-05, 
    3.066671e-05, 3.066652e-05, 3.066682e-05, 3.066672e-05, 3.066666e-05, 
    3.066669e-05, 3.066655e-05, 3.066652e-05, 3.066638e-05, 3.066645e-05, 
    3.066604e-05, 3.066622e-05, 3.066571e-05, 3.066585e-05, 3.066682e-05, 
    3.066677e-05, 3.066661e-05, 3.066668e-05, 3.066647e-05, 3.066642e-05, 
    3.066638e-05, 3.066632e-05, 3.066632e-05, 3.066628e-05, 3.066634e-05, 
    3.066628e-05, 3.066648e-05, 3.066639e-05, 3.066663e-05, 3.066657e-05, 
    3.06666e-05, 3.066663e-05, 3.066654e-05, 3.066644e-05, 3.066644e-05, 
    3.066641e-05, 3.066632e-05, 3.066647e-05, 3.066601e-05, 3.06663e-05, 
    3.066672e-05, 3.066663e-05, 3.066662e-05, 3.066665e-05, 3.066642e-05, 
    3.066651e-05, 3.066628e-05, 3.066634e-05, 3.066624e-05, 3.06663e-05, 
    3.06663e-05, 3.066636e-05, 3.06664e-05, 3.06665e-05, 3.066658e-05, 
    3.066665e-05, 3.066663e-05, 3.066656e-05, 3.066644e-05, 3.066631e-05, 
    3.066634e-05, 3.066625e-05, 3.066649e-05, 3.066639e-05, 3.066643e-05, 
    3.066633e-05, 3.066655e-05, 3.066636e-05, 3.066659e-05, 3.066657e-05, 
    3.066651e-05, 3.066638e-05, 3.066635e-05, 3.066632e-05, 3.066634e-05, 
    3.066643e-05, 3.066645e-05, 3.066651e-05, 3.066653e-05, 3.066658e-05, 
    3.066662e-05, 3.066658e-05, 3.066654e-05, 3.066643e-05, 3.066634e-05, 
    3.066623e-05, 3.06662e-05, 3.066608e-05, 3.066618e-05, 3.066601e-05, 
    3.066615e-05, 3.066591e-05, 3.066635e-05, 3.066616e-05, 3.066651e-05, 
    3.066647e-05, 3.06664e-05, 3.066624e-05, 3.066633e-05, 3.066623e-05, 
    3.066645e-05, 3.066656e-05, 3.066659e-05, 3.066664e-05, 3.066659e-05, 
    3.066659e-05, 3.066654e-05, 3.066656e-05, 3.066643e-05, 3.06665e-05, 
    3.06663e-05, 3.066623e-05, 3.066603e-05, 3.066591e-05, 3.066578e-05, 
    3.066573e-05, 3.066571e-05, 3.06657e-05 ;

 LITR1C_TO_SOIL1C =
  6.62691e-13, 6.643762e-13, 6.640488e-13, 6.654066e-13, 6.646538e-13, 
    6.655425e-13, 6.630331e-13, 6.644428e-13, 6.635432e-13, 6.628432e-13, 
    6.680372e-13, 6.654672e-13, 6.707045e-13, 6.690686e-13, 6.731752e-13, 
    6.704497e-13, 6.737243e-13, 6.730973e-13, 6.749849e-13, 6.744444e-13, 
    6.768547e-13, 6.752343e-13, 6.781035e-13, 6.764683e-13, 6.76724e-13, 
    6.751807e-13, 6.659854e-13, 6.677173e-13, 6.658826e-13, 6.661297e-13, 
    6.660189e-13, 6.646692e-13, 6.639881e-13, 6.625626e-13, 6.628216e-13, 
    6.638688e-13, 6.662408e-13, 6.654365e-13, 6.67464e-13, 6.674183e-13, 
    6.696719e-13, 6.686563e-13, 6.724392e-13, 6.713652e-13, 6.74467e-13, 
    6.736875e-13, 6.744303e-13, 6.742052e-13, 6.744333e-13, 6.732899e-13, 
    6.737798e-13, 6.727735e-13, 6.688464e-13, 6.700015e-13, 6.665534e-13, 
    6.644753e-13, 6.630949e-13, 6.62114e-13, 6.622528e-13, 6.62517e-13, 
    6.638749e-13, 6.65151e-13, 6.661225e-13, 6.66772e-13, 6.674117e-13, 
    6.693448e-13, 6.703682e-13, 6.72656e-13, 6.722439e-13, 6.729423e-13, 
    6.7361e-13, 6.747294e-13, 6.745453e-13, 6.750382e-13, 6.729243e-13, 
    6.743294e-13, 6.72009e-13, 6.72644e-13, 6.675835e-13, 6.656536e-13, 
    6.648308e-13, 6.641117e-13, 6.623593e-13, 6.635696e-13, 6.630926e-13, 
    6.642276e-13, 6.649481e-13, 6.645919e-13, 6.667898e-13, 6.659356e-13, 
    6.704288e-13, 6.684952e-13, 6.735321e-13, 6.723286e-13, 6.738205e-13, 
    6.730595e-13, 6.74363e-13, 6.7319e-13, 6.752218e-13, 6.756635e-13, 
    6.753616e-13, 6.765218e-13, 6.731248e-13, 6.744301e-13, 6.645818e-13, 
    6.646399e-13, 6.649107e-13, 6.637198e-13, 6.63647e-13, 6.625554e-13, 
    6.63527e-13, 6.639403e-13, 6.6499e-13, 6.656102e-13, 6.661996e-13, 
    6.674948e-13, 6.689395e-13, 6.70958e-13, 6.724066e-13, 6.733767e-13, 
    6.72782e-13, 6.73307e-13, 6.727201e-13, 6.72445e-13, 6.754979e-13, 
    6.737843e-13, 6.76355e-13, 6.762129e-13, 6.750499e-13, 6.762289e-13, 
    6.646807e-13, 6.643463e-13, 6.631842e-13, 6.640937e-13, 6.624365e-13, 
    6.633641e-13, 6.638971e-13, 6.65953e-13, 6.664048e-13, 6.66823e-13, 
    6.67649e-13, 6.687083e-13, 6.705643e-13, 6.721775e-13, 6.736489e-13, 
    6.735412e-13, 6.735791e-13, 6.739074e-13, 6.730937e-13, 6.740409e-13, 
    6.741996e-13, 6.737843e-13, 6.761939e-13, 6.755059e-13, 6.762099e-13, 
    6.757621e-13, 6.644551e-13, 6.650177e-13, 6.647137e-13, 6.652853e-13, 
    6.648824e-13, 6.666721e-13, 6.672083e-13, 6.69715e-13, 6.686873e-13, 
    6.703231e-13, 6.688537e-13, 6.691141e-13, 6.703756e-13, 6.689333e-13, 
    6.720882e-13, 6.699493e-13, 6.739201e-13, 6.717861e-13, 6.740537e-13, 
    6.736425e-13, 6.743234e-13, 6.749327e-13, 6.756993e-13, 6.771119e-13, 
    6.76785e-13, 6.779659e-13, 6.658563e-13, 6.665852e-13, 6.665214e-13, 
    6.67284e-13, 6.678478e-13, 6.690692e-13, 6.710257e-13, 6.702905e-13, 
    6.716405e-13, 6.719112e-13, 6.698603e-13, 6.711195e-13, 6.670731e-13, 
    6.677272e-13, 6.67338e-13, 6.659136e-13, 6.704594e-13, 6.68128e-13, 
    6.724304e-13, 6.711698e-13, 6.748458e-13, 6.730185e-13, 6.766049e-13, 
    6.781342e-13, 6.795737e-13, 6.812518e-13, 6.669832e-13, 6.664881e-13, 
    6.673748e-13, 6.686001e-13, 6.697371e-13, 6.712466e-13, 6.714012e-13, 
    6.716837e-13, 6.724156e-13, 6.730305e-13, 6.717726e-13, 6.731846e-13, 
    6.678781e-13, 6.706618e-13, 6.663005e-13, 6.676147e-13, 6.685281e-13, 
    6.681278e-13, 6.702065e-13, 6.706959e-13, 6.726825e-13, 6.71656e-13, 
    6.777566e-13, 6.750609e-13, 6.825293e-13, 6.804463e-13, 6.66315e-13, 
    6.669817e-13, 6.692991e-13, 6.68197e-13, 6.713476e-13, 6.721218e-13, 
    6.727512e-13, 6.735548e-13, 6.736418e-13, 6.741177e-13, 6.733377e-13, 
    6.74087e-13, 6.712498e-13, 6.725185e-13, 6.690349e-13, 6.698834e-13, 
    6.694932e-13, 6.690648e-13, 6.703864e-13, 6.717923e-13, 6.71823e-13, 
    6.722734e-13, 6.735407e-13, 6.713603e-13, 6.781029e-13, 6.739418e-13, 
    6.677083e-13, 6.689901e-13, 6.691739e-13, 6.686774e-13, 6.720442e-13, 
    6.708252e-13, 6.741062e-13, 6.732203e-13, 6.746716e-13, 6.739506e-13, 
    6.738444e-13, 6.729179e-13, 6.723405e-13, 6.708809e-13, 6.696924e-13, 
    6.687495e-13, 6.689688e-13, 6.700044e-13, 6.718784e-13, 6.736494e-13, 
    6.732616e-13, 6.745614e-13, 6.711194e-13, 6.725634e-13, 6.720053e-13, 
    6.734603e-13, 6.702708e-13, 6.729853e-13, 6.695758e-13, 6.698752e-13, 
    6.708009e-13, 6.726608e-13, 6.730729e-13, 6.735116e-13, 6.732411e-13, 
    6.719261e-13, 6.717108e-13, 6.707786e-13, 6.705208e-13, 6.698101e-13, 
    6.692212e-13, 6.697591e-13, 6.703237e-13, 6.719269e-13, 6.733697e-13, 
    6.749413e-13, 6.753259e-13, 6.771577e-13, 6.756658e-13, 6.78126e-13, 
    6.760334e-13, 6.796543e-13, 6.731434e-13, 6.759731e-13, 6.708433e-13, 
    6.71397e-13, 6.723973e-13, 6.746901e-13, 6.734534e-13, 6.748999e-13, 
    6.717024e-13, 6.700398e-13, 6.696101e-13, 6.688068e-13, 6.696285e-13, 
    6.695617e-13, 6.703475e-13, 6.700951e-13, 6.719801e-13, 6.709679e-13, 
    6.738416e-13, 6.748886e-13, 6.77842e-13, 6.796488e-13, 6.814864e-13, 
    6.822966e-13, 6.825432e-13, 6.826462e-13 ;

 LITR1C_vr =
  0.001751121, 0.001751114, 0.001751116, 0.00175111, 0.001751113, 0.00175111, 
    0.00175112, 0.001751114, 0.001751118, 0.00175112, 0.0017511, 0.00175111, 
    0.00175109, 0.001751096, 0.00175108, 0.001751091, 0.001751078, 
    0.00175108, 0.001751073, 0.001751075, 0.001751066, 0.001751072, 
    0.001751061, 0.001751067, 0.001751066, 0.001751072, 0.001751108, 
    0.001751101, 0.001751108, 0.001751108, 0.001751108, 0.001751113, 
    0.001751116, 0.001751121, 0.00175112, 0.001751116, 0.001751107, 
    0.00175111, 0.001751102, 0.001751103, 0.001751094, 0.001751098, 
    0.001751083, 0.001751087, 0.001751075, 0.001751078, 0.001751075, 
    0.001751076, 0.001751075, 0.00175108, 0.001751078, 0.001751082, 
    0.001751097, 0.001751092, 0.001751106, 0.001751114, 0.001751119, 
    0.001751123, 0.001751123, 0.001751121, 0.001751116, 0.001751111, 
    0.001751108, 0.001751105, 0.001751103, 0.001751095, 0.001751091, 
    0.001751082, 0.001751084, 0.001751081, 0.001751078, 0.001751074, 
    0.001751075, 0.001751073, 0.001751081, 0.001751076, 0.001751085, 
    0.001751082, 0.001751102, 0.001751109, 0.001751113, 0.001751115, 
    0.001751122, 0.001751117, 0.001751119, 0.001751115, 0.001751112, 
    0.001751113, 0.001751105, 0.001751108, 0.001751091, 0.001751098, 
    0.001751079, 0.001751083, 0.001751078, 0.001751081, 0.001751075, 
    0.00175108, 0.001751072, 0.00175107, 0.001751072, 0.001751067, 
    0.00175108, 0.001751075, 0.001751113, 0.001751113, 0.001751112, 
    0.001751117, 0.001751117, 0.001751121, 0.001751118, 0.001751116, 
    0.001751112, 0.001751109, 0.001751107, 0.001751102, 0.001751097, 
    0.001751089, 0.001751083, 0.001751079, 0.001751082, 0.00175108, 
    0.001751082, 0.001751083, 0.001751071, 0.001751078, 0.001751068, 
    0.001751068, 0.001751073, 0.001751068, 0.001751113, 0.001751114, 
    0.001751119, 0.001751115, 0.001751122, 0.001751118, 0.001751116, 
    0.001751108, 0.001751106, 0.001751105, 0.001751102, 0.001751098, 
    0.00175109, 0.001751084, 0.001751078, 0.001751079, 0.001751079, 
    0.001751077, 0.00175108, 0.001751077, 0.001751076, 0.001751078, 
    0.001751068, 0.001751071, 0.001751068, 0.00175107, 0.001751114, 
    0.001751112, 0.001751113, 0.001751111, 0.001751112, 0.001751105, 
    0.001751103, 0.001751094, 0.001751098, 0.001751091, 0.001751097, 
    0.001751096, 0.001751091, 0.001751097, 0.001751084, 0.001751093, 
    0.001751077, 0.001751086, 0.001751077, 0.001751078, 0.001751076, 
    0.001751073, 0.00175107, 0.001751065, 0.001751066, 0.001751062, 
    0.001751109, 0.001751106, 0.001751106, 0.001751103, 0.001751101, 
    0.001751096, 0.001751088, 0.001751091, 0.001751086, 0.001751085, 
    0.001751093, 0.001751088, 0.001751104, 0.001751101, 0.001751103, 
    0.001751108, 0.001751091, 0.0017511, 0.001751083, 0.001751088, 
    0.001751074, 0.001751081, 0.001751067, 0.001751061, 0.001751055, 
    0.001751049, 0.001751104, 0.001751106, 0.001751103, 0.001751098, 
    0.001751093, 0.001751088, 0.001751087, 0.001751086, 0.001751083, 
    0.001751081, 0.001751086, 0.00175108, 0.001751101, 0.00175109, 
    0.001751107, 0.001751102, 0.001751098, 0.0017511, 0.001751092, 
    0.00175109, 0.001751082, 0.001751086, 0.001751062, 0.001751073, 
    0.001751044, 0.001751052, 0.001751107, 0.001751104, 0.001751095, 
    0.001751099, 0.001751087, 0.001751084, 0.001751082, 0.001751079, 
    0.001751078, 0.001751076, 0.001751079, 0.001751077, 0.001751088, 
    0.001751083, 0.001751096, 0.001751093, 0.001751094, 0.001751096, 
    0.001751091, 0.001751086, 0.001751085, 0.001751084, 0.001751079, 
    0.001751087, 0.001751061, 0.001751077, 0.001751101, 0.001751096, 
    0.001751096, 0.001751098, 0.001751084, 0.001751089, 0.001751076, 
    0.00175108, 0.001751074, 0.001751077, 0.001751077, 0.001751081, 
    0.001751083, 0.001751089, 0.001751094, 0.001751097, 0.001751096, 
    0.001751092, 0.001751085, 0.001751078, 0.00175108, 0.001751075, 
    0.001751088, 0.001751082, 0.001751085, 0.001751079, 0.001751091, 
    0.001751081, 0.001751094, 0.001751093, 0.001751089, 0.001751082, 
    0.001751081, 0.001751079, 0.00175108, 0.001751085, 0.001751086, 
    0.001751089, 0.00175109, 0.001751093, 0.001751095, 0.001751093, 
    0.001751091, 0.001751085, 0.001751079, 0.001751073, 0.001751072, 
    0.001751065, 0.00175107, 0.001751061, 0.001751069, 0.001751055, 
    0.00175108, 0.001751069, 0.001751089, 0.001751087, 0.001751083, 
    0.001751074, 0.001751079, 0.001751073, 0.001751086, 0.001751092, 
    0.001751094, 0.001751097, 0.001751094, 0.001751094, 0.001751091, 
    0.001751092, 0.001751085, 0.001751089, 0.001751077, 0.001751073, 
    0.001751062, 0.001751055, 0.001751048, 0.001751045, 0.001751044, 
    0.001751043,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.732586e-07, 9.732549e-07, 9.732556e-07, 9.732527e-07, 9.732544e-07, 
    9.732524e-07, 9.732578e-07, 9.732548e-07, 9.732568e-07, 9.732582e-07, 
    9.73247e-07, 9.732526e-07, 9.732413e-07, 9.732448e-07, 9.73236e-07, 
    9.732419e-07, 9.732347e-07, 9.732361e-07, 9.73232e-07, 9.732332e-07, 
    9.73228e-07, 9.732315e-07, 9.732253e-07, 9.732288e-07, 9.732282e-07, 
    9.732316e-07, 9.732514e-07, 9.732478e-07, 9.732516e-07, 9.732512e-07, 
    9.732514e-07, 9.732543e-07, 9.732557e-07, 9.732588e-07, 9.732582e-07, 
    9.732561e-07, 9.73251e-07, 9.732527e-07, 9.732482e-07, 9.732483e-07, 
    9.732435e-07, 9.732457e-07, 9.732375e-07, 9.732398e-07, 9.732331e-07, 
    9.732348e-07, 9.732332e-07, 9.732337e-07, 9.732332e-07, 9.732357e-07, 
    9.732346e-07, 9.732368e-07, 9.732453e-07, 9.732428e-07, 9.732503e-07, 
    9.732547e-07, 9.732577e-07, 9.732598e-07, 9.732595e-07, 9.732589e-07, 
    9.73256e-07, 9.732532e-07, 9.732512e-07, 9.732497e-07, 9.732483e-07, 
    9.732443e-07, 9.73242e-07, 9.732371e-07, 9.73238e-07, 9.732364e-07, 
    9.73235e-07, 9.732325e-07, 9.73233e-07, 9.732319e-07, 9.732365e-07, 
    9.732335e-07, 9.732385e-07, 9.732371e-07, 9.73248e-07, 9.732522e-07, 
    9.732539e-07, 9.732555e-07, 9.732593e-07, 9.732566e-07, 9.732577e-07, 
    9.732553e-07, 9.732537e-07, 9.732545e-07, 9.732497e-07, 9.732515e-07, 
    9.732419e-07, 9.732461e-07, 9.732352e-07, 9.732378e-07, 9.732346e-07, 
    9.732362e-07, 9.732333e-07, 9.73236e-07, 9.732315e-07, 9.732306e-07, 
    9.732312e-07, 9.732287e-07, 9.732361e-07, 9.732332e-07, 9.732545e-07, 
    9.732544e-07, 9.732538e-07, 9.732563e-07, 9.732565e-07, 9.732589e-07, 
    9.732568e-07, 9.732559e-07, 9.732536e-07, 9.732523e-07, 9.73251e-07, 
    9.732482e-07, 9.732451e-07, 9.732407e-07, 9.732375e-07, 9.732355e-07, 
    9.732368e-07, 9.732356e-07, 9.732369e-07, 9.732375e-07, 9.73231e-07, 
    9.732346e-07, 9.73229e-07, 9.732294e-07, 9.732319e-07, 9.732294e-07, 
    9.732543e-07, 9.732551e-07, 9.732576e-07, 9.732555e-07, 9.732591e-07, 
    9.732571e-07, 9.73256e-07, 9.732515e-07, 9.732505e-07, 9.732496e-07, 
    9.732479e-07, 9.732456e-07, 9.732415e-07, 9.732381e-07, 9.732349e-07, 
    9.732352e-07, 9.73235e-07, 9.732344e-07, 9.732361e-07, 9.73234e-07, 
    9.732337e-07, 9.732346e-07, 9.732294e-07, 9.73231e-07, 9.732294e-07, 
    9.732304e-07, 9.732547e-07, 9.732536e-07, 9.732543e-07, 9.73253e-07, 
    9.732538e-07, 9.732499e-07, 9.732488e-07, 9.732435e-07, 9.732456e-07, 
    9.732421e-07, 9.732453e-07, 9.732447e-07, 9.73242e-07, 9.732451e-07, 
    9.732382e-07, 9.732429e-07, 9.732344e-07, 9.732389e-07, 9.73234e-07, 
    9.732349e-07, 9.732335e-07, 9.732321e-07, 9.732305e-07, 9.732274e-07, 
    9.732281e-07, 9.732256e-07, 9.732518e-07, 9.732502e-07, 9.732503e-07, 
    9.732487e-07, 9.732474e-07, 9.732448e-07, 9.732406e-07, 9.732422e-07, 
    9.732393e-07, 9.732387e-07, 9.732431e-07, 9.732404e-07, 9.732491e-07, 
    9.732477e-07, 9.732486e-07, 9.732516e-07, 9.732418e-07, 9.732469e-07, 
    9.732375e-07, 9.732403e-07, 9.732323e-07, 9.732363e-07, 9.732286e-07, 
    9.732253e-07, 9.732221e-07, 9.732184e-07, 9.732493e-07, 9.732504e-07, 
    9.732485e-07, 9.732458e-07, 9.732433e-07, 9.7324e-07, 9.732398e-07, 
    9.732391e-07, 9.732375e-07, 9.732363e-07, 9.732389e-07, 9.73236e-07, 
    9.732473e-07, 9.732414e-07, 9.732507e-07, 9.732479e-07, 9.73246e-07, 
    9.732469e-07, 9.732423e-07, 9.732413e-07, 9.73237e-07, 9.732393e-07, 
    9.732261e-07, 9.732319e-07, 9.732157e-07, 9.732203e-07, 9.732507e-07, 
    9.732493e-07, 9.732443e-07, 9.732466e-07, 9.732399e-07, 9.732382e-07, 
    9.732369e-07, 9.732352e-07, 9.732349e-07, 9.732339e-07, 9.732356e-07, 
    9.73234e-07, 9.7324e-07, 9.732373e-07, 9.732448e-07, 9.73243e-07, 
    9.732439e-07, 9.732448e-07, 9.73242e-07, 9.732389e-07, 9.732389e-07, 
    9.732379e-07, 9.732352e-07, 9.732398e-07, 9.732253e-07, 9.732343e-07, 
    9.732478e-07, 9.732449e-07, 9.732446e-07, 9.732456e-07, 9.732383e-07, 
    9.73241e-07, 9.732339e-07, 9.732358e-07, 9.732327e-07, 9.732343e-07, 
    9.732345e-07, 9.732365e-07, 9.732378e-07, 9.732408e-07, 9.732435e-07, 
    9.732455e-07, 9.732451e-07, 9.732428e-07, 9.732387e-07, 9.732349e-07, 
    9.732357e-07, 9.732329e-07, 9.732404e-07, 9.732372e-07, 9.732385e-07, 
    9.732353e-07, 9.732422e-07, 9.732363e-07, 9.732437e-07, 9.732431e-07, 
    9.732411e-07, 9.732371e-07, 9.732362e-07, 9.732352e-07, 9.732358e-07, 
    9.732387e-07, 9.732391e-07, 9.732411e-07, 9.732416e-07, 9.732432e-07, 
    9.732445e-07, 9.732433e-07, 9.732421e-07, 9.732387e-07, 9.732355e-07, 
    9.732321e-07, 9.732313e-07, 9.732273e-07, 9.732306e-07, 9.732253e-07, 
    9.732298e-07, 9.73222e-07, 9.73236e-07, 9.732299e-07, 9.73241e-07, 
    9.732398e-07, 9.732377e-07, 9.732327e-07, 9.732354e-07, 9.732322e-07, 
    9.732391e-07, 9.732427e-07, 9.732437e-07, 9.732454e-07, 9.732436e-07, 
    9.732437e-07, 9.732421e-07, 9.732425e-07, 9.732386e-07, 9.732407e-07, 
    9.732345e-07, 9.732322e-07, 9.732258e-07, 9.73222e-07, 9.73218e-07, 
    9.732163e-07, 9.732157e-07, 9.732155e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  -1.911706e-25, -2.058761e-25, -1.960724e-25, 1.088202e-24, -8.333079e-26, 
    -2.450906e-25, 8.333079e-25, 4.705739e-25, 8.137007e-25, -2.156797e-25, 
    -4.509666e-25, 3.039123e-25, 6.568427e-25, 6.568427e-25, 9.803622e-27, 
    -1.093104e-24, -8.137007e-25, 7.058608e-25, -2.450906e-25, 2.843051e-25, 
    9.803622e-27, 9.803622e-26, -8.333079e-26, -6.715481e-25, 7.450753e-25, 
    1.02938e-24, -6.274318e-25, -2.156797e-25, 3.088141e-25, -4.901811e-25, 
    1.127417e-25, -9.411477e-25, 6.960572e-25, 1.372507e-25, 2.107779e-25, 
    -2.941087e-26, 3.431268e-26, -3.333231e-25, 4.019485e-25, 6.47039e-25, 
    5.048866e-25, 6.764499e-25, -6.862535e-25, 8.284061e-25, 2.450905e-26, 
    -4.019485e-25, -3.872431e-25, 3.431268e-26, 4.313593e-25, -1.176435e-25, 
    3.235195e-25, -1.666616e-25, -2.745014e-25, -9.313441e-26, 4.215557e-25, 
    -5.588064e-25, -1.372507e-25, 4.901811e-25, -4.901811e-26, 2.205815e-25, 
    4.901811e-26, 7.107626e-25, -6.372354e-26, 7.842898e-26, -3.333231e-25, 
    2.941087e-26, 9.803622e-27, 2.156797e-25, 3.431268e-26, -4.901811e-26, 
    5.882173e-26, -3.823413e-25, -2.695996e-25, 3.529304e-25, 4.509666e-25, 
    5.784137e-25, -5.588064e-25, -2.548942e-25, -3.039123e-25, 4.166539e-25, 
    4.852793e-25, -2.548942e-25, 4.313593e-25, -3.137159e-25, -8.872278e-25, 
    3.921449e-26, 4.901811e-25, 2.794032e-25, 2.205815e-25, -1.441132e-24, 
    7.107626e-25, 1.421525e-25, 5.293956e-25, -3.480286e-25, -2.843051e-25, 
    3.676358e-25, 9.705585e-25, -6.274318e-25, 2.990105e-25, -3.333231e-25, 
    3.333231e-25, -9.803622e-27, -1.372507e-25, 1.81367e-25, 1.764652e-25, 
    -6.519409e-25, -4.754757e-25, 4.215557e-25, 7.891916e-25, 8.82326e-25, 
    2.548942e-25, 2.745014e-25, -3.333231e-25, -6.862535e-26, 6.274318e-25, 
    1.215649e-24, 2.646978e-25, 4.117521e-25, -4.65672e-25, 1.960724e-25, 
    -1.372507e-25, 5.19592e-25, 5.048866e-25, -2.450906e-25, 6.862535e-26, 
    4.901811e-26, -3.921449e-25, -1.078398e-25, 7.842898e-25, 3.725376e-25, 
    -1.764652e-25, -1.470543e-25, 4.313593e-25, -1.372507e-25, -9.313441e-26, 
    4.607703e-25, -1.911706e-25, 2.843051e-25, 2.646978e-25, 5.98021e-25, 
    3.431268e-25, -1.862688e-25, -8.82326e-26, 1.372507e-25, 2.646978e-25, 
    4.41163e-25, 9.803622e-27, 2.941087e-25, -6.862535e-25, -9.60755e-25, 
    6.078246e-25, 4.117521e-25, 5.882173e-26, 1.519561e-25, -4.999847e-25, 
    5.784137e-25, 7.646825e-25, 3.921449e-26, -8.137007e-25, 9.019333e-25, 
    -5.882173e-26, -1.81367e-25, 7.401734e-25, -3.137159e-25, -3.921449e-26, 
    4.901811e-27, -1.372507e-25, 5.097883e-25, 1.617598e-25, -1.274471e-25, 
    -3.186177e-25, 9.60755e-25, -1.176435e-25, -1.088202e-24, 4.019485e-25, 
    3.774394e-25, 5.882173e-26, 2.303851e-25, 8.431115e-25, 1.127417e-24, 
    1.02938e-25, 2.254833e-25, -7.842898e-25, 4.607703e-25, 9.803622e-27, 
    2.352869e-25, 3.137159e-25, 3.921449e-26, 1.960724e-25, 8.82326e-26, 
    -4.950829e-25, 4.803775e-25, 2.646978e-25, 4.901811e-27, 4.901811e-25, 
    1.862688e-25, 9.803622e-26, 1.666616e-25, 1.470543e-25, -1.56858e-25, 
    -2.843051e-25, 5.391992e-25, -1.02938e-25, 1.274471e-25, 6.421373e-25, 
    -2.695996e-25, 5.833155e-25, -3.137159e-25, 5.293956e-25, -2.941087e-26, 
    1.372507e-25, 7.842898e-26, -3.431268e-26, -2.548942e-25, -1.127417e-25, 
    8.529151e-25, 1.093104e-24, -3.235195e-25, 1.666616e-25, -1.960724e-25, 
    -7.401734e-25, -5.784137e-25, 6.617445e-25, 3.235195e-25, -4.901811e-26, 
    -2.892069e-25, -8.774241e-25, 5.391992e-25, 1.333293e-24, 2.156797e-25, 
    -6.862535e-26, 4.607703e-25, -5.490028e-25, -5.784137e-25, 4.901811e-26, 
    5.637083e-25, 4.264576e-25, -2.450906e-25, -2.058761e-25, 2.352869e-25, 
    1.56858e-25, 2.990105e-25, 2.843051e-25, -3.137159e-25, 4.803775e-25, 
    6.862535e-26, -7.842898e-26, 7.989952e-25, -3.284213e-25, 2.058761e-25, 
    -7.156644e-25, -4.901811e-26, 2.941087e-26, 6.862535e-25, 4.754757e-25, 
    -3.529304e-25, -4.068503e-25, -7.058608e-25, 4.607703e-25, -4.705739e-25, 
    2.59796e-25, 1.112711e-24, 3.970467e-25, -2.941087e-25, 6.862535e-26, 
    5.391992e-25, -1.372507e-25, -4.852793e-25, -2.695996e-25, -1.960724e-26, 
    -5.293956e-25, 7.940934e-25, 5.784137e-25, -5.882173e-26, -5.784137e-25, 
    -1.960724e-26, 8.82326e-26, -9.803622e-26, -7.646825e-25, 1.764652e-25, 
    5.588064e-25, 4.509666e-25, -3.529304e-25, -9.901658e-25, -2.941087e-26, 
    6.519409e-25, -4.362612e-25, -4.901811e-26, -2.156797e-25, -1.764652e-25, 
    -3.480286e-25, -1.862688e-25, -4.754757e-25, 5.98021e-25, -1.019577e-24, 
    4.313593e-25, 6.960572e-25, 1.078398e-24, -2.156797e-25, 2.646978e-25, 
    -3.872431e-25, -2.794032e-25, 1.666616e-25, 8.872278e-25, -1.176435e-25, 
    1.617598e-25, -2.450906e-25, 1.715634e-25, -2.352869e-25, -1.960724e-25, 
    6.715481e-25, 3.284213e-25, -1.666616e-25, 3.529304e-25, -6.862535e-26, 
    6.078246e-25, -1.274471e-25, 2.941087e-26, 2.941087e-25, -3.333231e-25, 
    -3.823413e-25, 7.842898e-26, 2.843051e-25, 3.62734e-25, 2.695996e-25, 
    6.078246e-25, 2.941087e-25, -2.646978e-25, 4.019485e-25, 6.372354e-25, 
    5.097883e-25, 3.137159e-25, 4.509666e-25, 6.176282e-25, -4.901811e-26, 
    -1.764652e-25, 1.02938e-24, 9.019333e-25,
  9.436424e-32, 9.436388e-32, 9.436395e-32, 9.436365e-32, 9.436381e-32, 
    9.436362e-32, 9.436417e-32, 9.436386e-32, 9.436406e-32, 9.436421e-32, 
    9.436308e-32, 9.436364e-32, 9.43625e-32, 9.436286e-32, 9.436197e-32, 
    9.436256e-32, 9.436185e-32, 9.436199e-32, 9.436157e-32, 9.436169e-32, 
    9.436117e-32, 9.436152e-32, 9.43609e-32, 9.436125e-32, 9.43612e-32, 
    9.436153e-32, 9.436353e-32, 9.436315e-32, 9.436355e-32, 9.43635e-32, 
    9.436352e-32, 9.436381e-32, 9.436396e-32, 9.436427e-32, 9.436421e-32, 
    9.436398e-32, 9.436347e-32, 9.436364e-32, 9.436321e-32, 9.436321e-32, 
    9.436273e-32, 9.436295e-32, 9.436213e-32, 9.436236e-32, 9.436169e-32, 
    9.436186e-32, 9.436169e-32, 9.436175e-32, 9.436169e-32, 9.436195e-32, 
    9.436183e-32, 9.436206e-32, 9.436291e-32, 9.436266e-32, 9.43634e-32, 
    9.436386e-32, 9.436415e-32, 9.436437e-32, 9.436434e-32, 9.436428e-32, 
    9.436398e-32, 9.436371e-32, 9.43635e-32, 9.436336e-32, 9.436321e-32, 
    9.43628e-32, 9.436257e-32, 9.436208e-32, 9.436217e-32, 9.436202e-32, 
    9.436187e-32, 9.436163e-32, 9.436167e-32, 9.436156e-32, 9.436202e-32, 
    9.436172e-32, 9.436222e-32, 9.436208e-32, 9.436318e-32, 9.43636e-32, 
    9.436378e-32, 9.436393e-32, 9.436431e-32, 9.436405e-32, 9.436415e-32, 
    9.436391e-32, 9.436375e-32, 9.436383e-32, 9.436335e-32, 9.436354e-32, 
    9.436256e-32, 9.436299e-32, 9.436189e-32, 9.436215e-32, 9.436183e-32, 
    9.436199e-32, 9.436171e-32, 9.436196e-32, 9.436152e-32, 9.436143e-32, 
    9.436149e-32, 9.436124e-32, 9.436198e-32, 9.436169e-32, 9.436383e-32, 
    9.436382e-32, 9.436376e-32, 9.436402e-32, 9.436403e-32, 9.436427e-32, 
    9.436406e-32, 9.436397e-32, 9.436374e-32, 9.436361e-32, 9.436348e-32, 
    9.43632e-32, 9.436289e-32, 9.436245e-32, 9.436213e-32, 9.436192e-32, 
    9.436205e-32, 9.436194e-32, 9.436207e-32, 9.436213e-32, 9.436146e-32, 
    9.436183e-32, 9.436127e-32, 9.436131e-32, 9.436156e-32, 9.43613e-32, 
    9.436381e-32, 9.436388e-32, 9.436414e-32, 9.436394e-32, 9.43643e-32, 
    9.43641e-32, 9.436398e-32, 9.436353e-32, 9.436344e-32, 9.436334e-32, 
    9.436317e-32, 9.436294e-32, 9.436253e-32, 9.436219e-32, 9.436186e-32, 
    9.436189e-32, 9.436188e-32, 9.436181e-32, 9.436199e-32, 9.436178e-32, 
    9.436175e-32, 9.436183e-32, 9.436131e-32, 9.436146e-32, 9.436131e-32, 
    9.43614e-32, 9.436386e-32, 9.436374e-32, 9.43638e-32, 9.436368e-32, 
    9.436377e-32, 9.436338e-32, 9.436326e-32, 9.436271e-32, 9.436294e-32, 
    9.436259e-32, 9.43629e-32, 9.436285e-32, 9.436257e-32, 9.436289e-32, 
    9.43622e-32, 9.436267e-32, 9.43618e-32, 9.436227e-32, 9.436177e-32, 
    9.436187e-32, 9.436172e-32, 9.436159e-32, 9.436142e-32, 9.436111e-32, 
    9.436119e-32, 9.436093e-32, 9.436356e-32, 9.43634e-32, 9.436341e-32, 
    9.436324e-32, 9.436312e-32, 9.436286e-32, 9.436243e-32, 9.436259e-32, 
    9.43623e-32, 9.436224e-32, 9.436269e-32, 9.436242e-32, 9.436329e-32, 
    9.436315e-32, 9.436323e-32, 9.436354e-32, 9.436256e-32, 9.436306e-32, 
    9.436213e-32, 9.43624e-32, 9.43616e-32, 9.4362e-32, 9.436122e-32, 
    9.436089e-32, 9.436058e-32, 9.436022e-32, 9.436331e-32, 9.436342e-32, 
    9.436323e-32, 9.436296e-32, 9.436271e-32, 9.436239e-32, 9.436235e-32, 
    9.436229e-32, 9.436213e-32, 9.4362e-32, 9.436227e-32, 9.436196e-32, 
    9.436311e-32, 9.436252e-32, 9.436346e-32, 9.436317e-32, 9.436297e-32, 
    9.436306e-32, 9.436261e-32, 9.43625e-32, 9.436207e-32, 9.43623e-32, 
    9.436098e-32, 9.436156e-32, 9.435993e-32, 9.436039e-32, 9.436346e-32, 
    9.436331e-32, 9.436281e-32, 9.436305e-32, 9.436236e-32, 9.43622e-32, 
    9.436206e-32, 9.436189e-32, 9.436187e-32, 9.436176e-32, 9.436193e-32, 
    9.436177e-32, 9.436239e-32, 9.436211e-32, 9.436287e-32, 9.436268e-32, 
    9.436277e-32, 9.436286e-32, 9.436257e-32, 9.436227e-32, 9.436226e-32, 
    9.436216e-32, 9.436189e-32, 9.436236e-32, 9.43609e-32, 9.43618e-32, 
    9.436316e-32, 9.436287e-32, 9.436283e-32, 9.436294e-32, 9.436222e-32, 
    9.436248e-32, 9.436176e-32, 9.436196e-32, 9.436165e-32, 9.43618e-32, 
    9.436182e-32, 9.436202e-32, 9.436215e-32, 9.436246e-32, 9.436272e-32, 
    9.436293e-32, 9.436288e-32, 9.436266e-32, 9.436225e-32, 9.436186e-32, 
    9.436195e-32, 9.436167e-32, 9.436242e-32, 9.43621e-32, 9.436222e-32, 
    9.43619e-32, 9.43626e-32, 9.436201e-32, 9.436275e-32, 9.436269e-32, 
    9.436248e-32, 9.436208e-32, 9.436199e-32, 9.436189e-32, 9.436195e-32, 
    9.436224e-32, 9.436229e-32, 9.436249e-32, 9.436254e-32, 9.43627e-32, 
    9.436283e-32, 9.436271e-32, 9.436259e-32, 9.436224e-32, 9.436193e-32, 
    9.436159e-32, 9.43615e-32, 9.43611e-32, 9.436143e-32, 9.436089e-32, 
    9.436135e-32, 9.436056e-32, 9.436197e-32, 9.436136e-32, 9.436247e-32, 
    9.436235e-32, 9.436213e-32, 9.436164e-32, 9.436191e-32, 9.436159e-32, 
    9.436229e-32, 9.436265e-32, 9.436274e-32, 9.436291e-32, 9.436274e-32, 
    9.436275e-32, 9.436258e-32, 9.436263e-32, 9.436223e-32, 9.436244e-32, 
    9.436182e-32, 9.43616e-32, 9.436096e-32, 9.436056e-32, 9.436016e-32, 
    9.435999e-32, 9.435993e-32, 9.435991e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.673629e-14, 4.685513e-14, 4.683205e-14, 4.692781e-14, 4.687472e-14, 
    4.693739e-14, 4.676041e-14, 4.685983e-14, 4.679639e-14, 4.674702e-14, 
    4.711333e-14, 4.693208e-14, 4.730144e-14, 4.718606e-14, 4.747569e-14, 
    4.728347e-14, 4.751441e-14, 4.747019e-14, 4.760332e-14, 4.75652e-14, 
    4.773519e-14, 4.76209e-14, 4.782325e-14, 4.770793e-14, 4.772596e-14, 
    4.761713e-14, 4.696862e-14, 4.709077e-14, 4.696137e-14, 4.69788e-14, 
    4.697099e-14, 4.68758e-14, 4.682776e-14, 4.672723e-14, 4.67455e-14, 
    4.681935e-14, 4.698664e-14, 4.692991e-14, 4.70729e-14, 4.706968e-14, 
    4.722862e-14, 4.715699e-14, 4.742378e-14, 4.734804e-14, 4.756679e-14, 
    4.751182e-14, 4.75642e-14, 4.754833e-14, 4.756441e-14, 4.748377e-14, 
    4.751833e-14, 4.744735e-14, 4.71704e-14, 4.725186e-14, 4.700868e-14, 
    4.686212e-14, 4.676477e-14, 4.66956e-14, 4.670538e-14, 4.672401e-14, 
    4.681978e-14, 4.690978e-14, 4.69783e-14, 4.70241e-14, 4.706921e-14, 
    4.720555e-14, 4.727772e-14, 4.743907e-14, 4.741001e-14, 4.745926e-14, 
    4.750635e-14, 4.75853e-14, 4.757231e-14, 4.760707e-14, 4.745799e-14, 
    4.755708e-14, 4.739344e-14, 4.743822e-14, 4.708133e-14, 4.694522e-14, 
    4.688719e-14, 4.683648e-14, 4.671289e-14, 4.679825e-14, 4.676461e-14, 
    4.684466e-14, 4.689547e-14, 4.687035e-14, 4.702535e-14, 4.696511e-14, 
    4.7282e-14, 4.714563e-14, 4.750086e-14, 4.741598e-14, 4.75212e-14, 
    4.746753e-14, 4.755946e-14, 4.747673e-14, 4.762002e-14, 4.765118e-14, 
    4.762988e-14, 4.77117e-14, 4.747213e-14, 4.756419e-14, 4.686964e-14, 
    4.687373e-14, 4.689283e-14, 4.680884e-14, 4.680371e-14, 4.672672e-14, 
    4.679524e-14, 4.682439e-14, 4.689843e-14, 4.694216e-14, 4.698373e-14, 
    4.707507e-14, 4.717697e-14, 4.731931e-14, 4.742148e-14, 4.748989e-14, 
    4.744796e-14, 4.748498e-14, 4.744359e-14, 4.742419e-14, 4.763949e-14, 
    4.751864e-14, 4.769994e-14, 4.768992e-14, 4.760789e-14, 4.769105e-14, 
    4.687661e-14, 4.685303e-14, 4.677107e-14, 4.683522e-14, 4.671834e-14, 
    4.678376e-14, 4.682135e-14, 4.696634e-14, 4.69982e-14, 4.70277e-14, 
    4.708596e-14, 4.716065e-14, 4.729155e-14, 4.740532e-14, 4.750909e-14, 
    4.75015e-14, 4.750417e-14, 4.752732e-14, 4.746994e-14, 4.753674e-14, 
    4.754793e-14, 4.751864e-14, 4.768858e-14, 4.764006e-14, 4.768971e-14, 
    4.765813e-14, 4.68607e-14, 4.690038e-14, 4.687894e-14, 4.691925e-14, 
    4.689084e-14, 4.701706e-14, 4.705487e-14, 4.723165e-14, 4.715918e-14, 
    4.727454e-14, 4.717091e-14, 4.718927e-14, 4.727824e-14, 4.717652e-14, 
    4.739903e-14, 4.724818e-14, 4.752822e-14, 4.737772e-14, 4.753764e-14, 
    4.750864e-14, 4.755666e-14, 4.759964e-14, 4.76537e-14, 4.775332e-14, 
    4.773027e-14, 4.781355e-14, 4.695952e-14, 4.701092e-14, 4.700643e-14, 
    4.706021e-14, 4.709997e-14, 4.718611e-14, 4.73241e-14, 4.727224e-14, 
    4.736745e-14, 4.738654e-14, 4.72419e-14, 4.733071e-14, 4.704533e-14, 
    4.709146e-14, 4.706402e-14, 4.696356e-14, 4.728415e-14, 4.711973e-14, 
    4.742316e-14, 4.733425e-14, 4.759351e-14, 4.746463e-14, 4.771757e-14, 
    4.782542e-14, 4.792694e-14, 4.804529e-14, 4.7039e-14, 4.700408e-14, 
    4.706662e-14, 4.715303e-14, 4.723321e-14, 4.733967e-14, 4.735057e-14, 
    4.73705e-14, 4.742211e-14, 4.746548e-14, 4.737677e-14, 4.747635e-14, 
    4.710211e-14, 4.729842e-14, 4.699085e-14, 4.708353e-14, 4.714794e-14, 
    4.711972e-14, 4.726632e-14, 4.730083e-14, 4.744093e-14, 4.736855e-14, 
    4.779879e-14, 4.760867e-14, 4.813539e-14, 4.798848e-14, 4.699187e-14, 
    4.703889e-14, 4.720232e-14, 4.71246e-14, 4.734679e-14, 4.740139e-14, 
    4.744578e-14, 4.750245e-14, 4.750859e-14, 4.754215e-14, 4.748715e-14, 
    4.753999e-14, 4.73399e-14, 4.742937e-14, 4.718369e-14, 4.724353e-14, 
    4.721601e-14, 4.71858e-14, 4.727901e-14, 4.737816e-14, 4.738032e-14, 
    4.741208e-14, 4.750146e-14, 4.734769e-14, 4.782321e-14, 4.752975e-14, 
    4.709013e-14, 4.718053e-14, 4.719349e-14, 4.715848e-14, 4.739592e-14, 
    4.730995e-14, 4.754134e-14, 4.747887e-14, 4.758122e-14, 4.753037e-14, 
    4.752289e-14, 4.745754e-14, 4.741682e-14, 4.731388e-14, 4.723006e-14, 
    4.716356e-14, 4.717903e-14, 4.725206e-14, 4.738423e-14, 4.750913e-14, 
    4.748178e-14, 4.757345e-14, 4.73307e-14, 4.743254e-14, 4.739317e-14, 
    4.749579e-14, 4.727085e-14, 4.74623e-14, 4.722184e-14, 4.724296e-14, 
    4.730824e-14, 4.743941e-14, 4.746847e-14, 4.749942e-14, 4.748033e-14, 
    4.738759e-14, 4.737241e-14, 4.730666e-14, 4.728848e-14, 4.723836e-14, 
    4.719683e-14, 4.723477e-14, 4.727459e-14, 4.738765e-14, 4.74894e-14, 
    4.760024e-14, 4.762736e-14, 4.775655e-14, 4.765134e-14, 4.782484e-14, 
    4.767726e-14, 4.793263e-14, 4.747345e-14, 4.7673e-14, 4.731123e-14, 
    4.735028e-14, 4.742082e-14, 4.758252e-14, 4.749531e-14, 4.759732e-14, 
    4.737182e-14, 4.725456e-14, 4.722426e-14, 4.71676e-14, 4.722555e-14, 
    4.722084e-14, 4.727626e-14, 4.725846e-14, 4.73914e-14, 4.732001e-14, 
    4.752269e-14, 4.759653e-14, 4.780481e-14, 4.793223e-14, 4.806184e-14, 
    4.811897e-14, 4.813636e-14, 4.814362e-14 ;

 LITR1N_vr =
  5.557407e-05, 5.557386e-05, 5.55739e-05, 5.557374e-05, 5.557383e-05, 
    5.557372e-05, 5.557403e-05, 5.557386e-05, 5.557396e-05, 5.557405e-05, 
    5.557341e-05, 5.557373e-05, 5.557308e-05, 5.557328e-05, 5.557278e-05, 
    5.557311e-05, 5.557271e-05, 5.557279e-05, 5.557255e-05, 5.557262e-05, 
    5.557232e-05, 5.557252e-05, 5.557217e-05, 5.557237e-05, 5.557234e-05, 
    5.557253e-05, 5.557366e-05, 5.557345e-05, 5.557368e-05, 5.557365e-05, 
    5.557366e-05, 5.557383e-05, 5.557391e-05, 5.557408e-05, 5.557406e-05, 
    5.557392e-05, 5.557363e-05, 5.557373e-05, 5.557348e-05, 5.557349e-05, 
    5.557321e-05, 5.557333e-05, 5.557287e-05, 5.5573e-05, 5.557262e-05, 
    5.557271e-05, 5.557262e-05, 5.557265e-05, 5.557262e-05, 5.557276e-05, 
    5.55727e-05, 5.557283e-05, 5.557331e-05, 5.557317e-05, 5.557359e-05, 
    5.557385e-05, 5.557402e-05, 5.557414e-05, 5.557412e-05, 5.557409e-05, 
    5.557392e-05, 5.557377e-05, 5.557365e-05, 5.557357e-05, 5.557349e-05, 
    5.557325e-05, 5.557312e-05, 5.557284e-05, 5.557289e-05, 5.557281e-05, 
    5.557272e-05, 5.557259e-05, 5.557261e-05, 5.557255e-05, 5.557281e-05, 
    5.557264e-05, 5.557292e-05, 5.557284e-05, 5.557347e-05, 5.557371e-05, 
    5.557381e-05, 5.55739e-05, 5.557411e-05, 5.557396e-05, 5.557402e-05, 
    5.557388e-05, 5.557379e-05, 5.557384e-05, 5.557356e-05, 5.557367e-05, 
    5.557312e-05, 5.557335e-05, 5.557273e-05, 5.557288e-05, 5.55727e-05, 
    5.557279e-05, 5.557263e-05, 5.557277e-05, 5.557252e-05, 5.557247e-05, 
    5.557251e-05, 5.557236e-05, 5.557279e-05, 5.557262e-05, 5.557384e-05, 
    5.557383e-05, 5.55738e-05, 5.557394e-05, 5.557395e-05, 5.557409e-05, 
    5.557397e-05, 5.557392e-05, 5.557379e-05, 5.557371e-05, 5.557364e-05, 
    5.557348e-05, 5.55733e-05, 5.557305e-05, 5.557287e-05, 5.557275e-05, 
    5.557283e-05, 5.557276e-05, 5.557283e-05, 5.557287e-05, 5.557249e-05, 
    5.55727e-05, 5.557239e-05, 5.55724e-05, 5.557255e-05, 5.55724e-05, 
    5.557383e-05, 5.557387e-05, 5.557401e-05, 5.55739e-05, 5.55741e-05, 
    5.557399e-05, 5.557392e-05, 5.557367e-05, 5.557361e-05, 5.557356e-05, 
    5.557346e-05, 5.557333e-05, 5.55731e-05, 5.55729e-05, 5.557272e-05, 
    5.557273e-05, 5.557273e-05, 5.557269e-05, 5.557279e-05, 5.557267e-05, 
    5.557265e-05, 5.55727e-05, 5.55724e-05, 5.557249e-05, 5.55724e-05, 
    5.557246e-05, 5.557385e-05, 5.557378e-05, 5.557382e-05, 5.557375e-05, 
    5.55738e-05, 5.557358e-05, 5.557351e-05, 5.55732e-05, 5.557333e-05, 
    5.557313e-05, 5.557331e-05, 5.557328e-05, 5.557312e-05, 5.55733e-05, 
    5.557291e-05, 5.557317e-05, 5.557269e-05, 5.557295e-05, 5.557267e-05, 
    5.557272e-05, 5.557264e-05, 5.557256e-05, 5.557247e-05, 5.557229e-05, 
    5.557233e-05, 5.557219e-05, 5.557368e-05, 5.557359e-05, 5.55736e-05, 
    5.55735e-05, 5.557343e-05, 5.557328e-05, 5.557304e-05, 5.557313e-05, 
    5.557297e-05, 5.557293e-05, 5.557319e-05, 5.557303e-05, 5.557353e-05, 
    5.557345e-05, 5.55735e-05, 5.557367e-05, 5.557311e-05, 5.55734e-05, 
    5.557287e-05, 5.557303e-05, 5.557257e-05, 5.55728e-05, 5.557236e-05, 
    5.557217e-05, 5.557199e-05, 5.557178e-05, 5.557354e-05, 5.55736e-05, 
    5.557349e-05, 5.557334e-05, 5.55732e-05, 5.557301e-05, 5.5573e-05, 
    5.557296e-05, 5.557287e-05, 5.55728e-05, 5.557295e-05, 5.557277e-05, 
    5.557343e-05, 5.557309e-05, 5.557363e-05, 5.557346e-05, 5.557335e-05, 
    5.55734e-05, 5.557314e-05, 5.557308e-05, 5.557284e-05, 5.557296e-05, 
    5.557221e-05, 5.557255e-05, 5.557163e-05, 5.557188e-05, 5.557362e-05, 
    5.557354e-05, 5.557325e-05, 5.557339e-05, 5.5573e-05, 5.557291e-05, 
    5.557283e-05, 5.557273e-05, 5.557272e-05, 5.557266e-05, 5.557276e-05, 
    5.557267e-05, 5.557301e-05, 5.557286e-05, 5.557329e-05, 5.557318e-05, 
    5.557323e-05, 5.557328e-05, 5.557312e-05, 5.557295e-05, 5.557295e-05, 
    5.557289e-05, 5.557273e-05, 5.5573e-05, 5.557217e-05, 5.557268e-05, 
    5.557345e-05, 5.557329e-05, 5.557327e-05, 5.557333e-05, 5.557292e-05, 
    5.557307e-05, 5.557266e-05, 5.557277e-05, 5.557259e-05, 5.557268e-05, 
    5.557269e-05, 5.557281e-05, 5.557288e-05, 5.557306e-05, 5.557321e-05, 
    5.557332e-05, 5.557329e-05, 5.557317e-05, 5.557294e-05, 5.557272e-05, 
    5.557277e-05, 5.557261e-05, 5.557303e-05, 5.557285e-05, 5.557292e-05, 
    5.557274e-05, 5.557313e-05, 5.55728e-05, 5.557322e-05, 5.557319e-05, 
    5.557307e-05, 5.557284e-05, 5.557279e-05, 5.557273e-05, 5.557277e-05, 
    5.557293e-05, 5.557296e-05, 5.557307e-05, 5.557311e-05, 5.557319e-05, 
    5.557327e-05, 5.55732e-05, 5.557313e-05, 5.557293e-05, 5.557275e-05, 
    5.557256e-05, 5.557251e-05, 5.557229e-05, 5.557247e-05, 5.557217e-05, 
    5.557243e-05, 5.557198e-05, 5.557278e-05, 5.557243e-05, 5.557307e-05, 
    5.5573e-05, 5.557287e-05, 5.557259e-05, 5.557274e-05, 5.557256e-05, 
    5.557296e-05, 5.557316e-05, 5.557322e-05, 5.557332e-05, 5.557321e-05, 
    5.557322e-05, 5.557313e-05, 5.557316e-05, 5.557292e-05, 5.557305e-05, 
    5.557269e-05, 5.557257e-05, 5.55722e-05, 5.557198e-05, 5.557175e-05, 
    5.557165e-05, 5.557162e-05, 5.557161e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  8.099557e-13, 8.120153e-13, 8.116153e-13, 8.132747e-13, 8.123546e-13, 
    8.134408e-13, 8.103738e-13, 8.120967e-13, 8.109972e-13, 8.101417e-13, 
    8.164899e-13, 8.133488e-13, 8.197499e-13, 8.177505e-13, 8.227697e-13, 
    8.194385e-13, 8.234408e-13, 8.226744e-13, 8.249816e-13, 8.24321e-13, 
    8.272669e-13, 8.252864e-13, 8.287931e-13, 8.267946e-13, 8.27107e-13, 
    8.252209e-13, 8.139821e-13, 8.160989e-13, 8.138565e-13, 8.141585e-13, 
    8.140232e-13, 8.123734e-13, 8.11541e-13, 8.097987e-13, 8.101153e-13, 
    8.113951e-13, 8.142944e-13, 8.133112e-13, 8.157894e-13, 8.157335e-13, 
    8.184879e-13, 8.172465e-13, 8.218701e-13, 8.205575e-13, 8.243486e-13, 
    8.233959e-13, 8.243037e-13, 8.240286e-13, 8.243073e-13, 8.229098e-13, 
    8.235087e-13, 8.222787e-13, 8.17479e-13, 8.188907e-13, 8.146763e-13, 
    8.121364e-13, 8.104493e-13, 8.092505e-13, 8.0942e-13, 8.09743e-13, 
    8.114026e-13, 8.129623e-13, 8.141497e-13, 8.149435e-13, 8.157254e-13, 
    8.180881e-13, 8.193389e-13, 8.221351e-13, 8.216314e-13, 8.224851e-13, 
    8.233011e-13, 8.246693e-13, 8.244443e-13, 8.250467e-13, 8.22463e-13, 
    8.241804e-13, 8.213443e-13, 8.221204e-13, 8.159354e-13, 8.135766e-13, 
    8.125709e-13, 8.116921e-13, 8.095503e-13, 8.110295e-13, 8.104465e-13, 
    8.118337e-13, 8.127143e-13, 8.12279e-13, 8.149652e-13, 8.139213e-13, 
    8.19413e-13, 8.170497e-13, 8.232059e-13, 8.217349e-13, 8.235584e-13, 
    8.226283e-13, 8.242215e-13, 8.227877e-13, 8.25271e-13, 8.25811e-13, 
    8.25442e-13, 8.268599e-13, 8.227081e-13, 8.243035e-13, 8.122666e-13, 
    8.123377e-13, 8.126687e-13, 8.112131e-13, 8.111242e-13, 8.097899e-13, 
    8.109774e-13, 8.114826e-13, 8.127656e-13, 8.135236e-13, 8.14244e-13, 
    8.15827e-13, 8.175928e-13, 8.200597e-13, 8.218302e-13, 8.230159e-13, 
    8.222892e-13, 8.229308e-13, 8.222134e-13, 8.218772e-13, 8.256085e-13, 
    8.235141e-13, 8.266561e-13, 8.264824e-13, 8.250609e-13, 8.26502e-13, 
    8.123875e-13, 8.119788e-13, 8.105585e-13, 8.116701e-13, 8.096446e-13, 
    8.107784e-13, 8.114298e-13, 8.139426e-13, 8.144948e-13, 8.150059e-13, 
    8.160155e-13, 8.1731e-13, 8.195786e-13, 8.215503e-13, 8.233487e-13, 
    8.23217e-13, 8.232633e-13, 8.236645e-13, 8.226702e-13, 8.238278e-13, 
    8.240217e-13, 8.235142e-13, 8.264592e-13, 8.256184e-13, 8.264788e-13, 
    8.259314e-13, 8.121118e-13, 8.127994e-13, 8.124279e-13, 8.131264e-13, 
    8.126341e-13, 8.148215e-13, 8.154768e-13, 8.185405e-13, 8.172844e-13, 
    8.192838e-13, 8.174878e-13, 8.178061e-13, 8.19348e-13, 8.175851e-13, 
    8.214412e-13, 8.188269e-13, 8.236802e-13, 8.210719e-13, 8.238434e-13, 
    8.233409e-13, 8.241731e-13, 8.249178e-13, 8.258547e-13, 8.275812e-13, 
    8.271817e-13, 8.286249e-13, 8.138244e-13, 8.147152e-13, 8.146373e-13, 
    8.155694e-13, 8.162584e-13, 8.177513e-13, 8.201426e-13, 8.192439e-13, 
    8.208939e-13, 8.212248e-13, 8.187182e-13, 8.202572e-13, 8.153115e-13, 
    8.16111e-13, 8.156354e-13, 8.138944e-13, 8.194504e-13, 8.166009e-13, 
    8.218594e-13, 8.203186e-13, 8.248116e-13, 8.225782e-13, 8.269616e-13, 
    8.288307e-13, 8.3059e-13, 8.326411e-13, 8.152017e-13, 8.145966e-13, 
    8.156804e-13, 8.171779e-13, 8.185675e-13, 8.204125e-13, 8.206015e-13, 
    8.209467e-13, 8.218413e-13, 8.225928e-13, 8.210554e-13, 8.227812e-13, 
    8.162954e-13, 8.196977e-13, 8.143673e-13, 8.159735e-13, 8.170898e-13, 
    8.166007e-13, 8.191413e-13, 8.197394e-13, 8.221674e-13, 8.209129e-13, 
    8.283692e-13, 8.250744e-13, 8.342026e-13, 8.316565e-13, 8.14385e-13, 
    8.151998e-13, 8.180322e-13, 8.166853e-13, 8.205359e-13, 8.214822e-13, 
    8.222515e-13, 8.232336e-13, 8.2334e-13, 8.239216e-13, 8.229683e-13, 
    8.238841e-13, 8.204165e-13, 8.219671e-13, 8.177093e-13, 8.187463e-13, 
    8.182694e-13, 8.177459e-13, 8.193612e-13, 8.210795e-13, 8.21117e-13, 
    8.216674e-13, 8.232163e-13, 8.205515e-13, 8.287925e-13, 8.237066e-13, 
    8.160879e-13, 8.176546e-13, 8.178792e-13, 8.172724e-13, 8.213873e-13, 
    8.198974e-13, 8.239076e-13, 8.228248e-13, 8.245987e-13, 8.237174e-13, 
    8.235877e-13, 8.224552e-13, 8.217495e-13, 8.199656e-13, 8.185129e-13, 
    8.173605e-13, 8.176286e-13, 8.188943e-13, 8.211848e-13, 8.233493e-13, 
    8.228752e-13, 8.244639e-13, 8.202569e-13, 8.220219e-13, 8.213397e-13, 
    8.23118e-13, 8.192199e-13, 8.225376e-13, 8.183705e-13, 8.187364e-13, 
    8.198678e-13, 8.22141e-13, 8.226447e-13, 8.231809e-13, 8.228502e-13, 
    8.21243e-13, 8.209799e-13, 8.198405e-13, 8.195254e-13, 8.186568e-13, 
    8.17937e-13, 8.185945e-13, 8.192845e-13, 8.21244e-13, 8.230075e-13, 
    8.249283e-13, 8.253983e-13, 8.276372e-13, 8.258138e-13, 8.288206e-13, 
    8.26263e-13, 8.306886e-13, 8.227308e-13, 8.261893e-13, 8.199195e-13, 
    8.205963e-13, 8.218188e-13, 8.246212e-13, 8.231097e-13, 8.248777e-13, 
    8.209696e-13, 8.189376e-13, 8.184123e-13, 8.174304e-13, 8.184348e-13, 
    8.183531e-13, 8.193136e-13, 8.190051e-13, 8.21309e-13, 8.200719e-13, 
    8.235842e-13, 8.248639e-13, 8.284735e-13, 8.306818e-13, 8.329279e-13, 
    8.339181e-13, 8.342194e-13, 8.343453e-13 ;

 LITR2C =
  1.939584e-05, 1.939582e-05, 1.939582e-05, 1.939581e-05, 1.939581e-05, 
    1.93958e-05, 1.939583e-05, 1.939582e-05, 1.939583e-05, 1.939583e-05, 
    1.939578e-05, 1.939581e-05, 1.939575e-05, 1.939576e-05, 1.939572e-05, 
    1.939575e-05, 1.939571e-05, 1.939572e-05, 1.93957e-05, 1.93957e-05, 
    1.939568e-05, 1.939569e-05, 1.939566e-05, 1.939568e-05, 1.939568e-05, 
    1.939569e-05, 1.93958e-05, 1.939578e-05, 1.93958e-05, 1.93958e-05, 
    1.93958e-05, 1.939581e-05, 1.939582e-05, 1.939584e-05, 1.939583e-05, 
    1.939582e-05, 1.93958e-05, 1.939581e-05, 1.939578e-05, 1.939578e-05, 
    1.939576e-05, 1.939577e-05, 1.939573e-05, 1.939574e-05, 1.93957e-05, 
    1.939571e-05, 1.93957e-05, 1.939571e-05, 1.93957e-05, 1.939572e-05, 
    1.939571e-05, 1.939572e-05, 1.939577e-05, 1.939575e-05, 1.939579e-05, 
    1.939582e-05, 1.939583e-05, 1.939584e-05, 1.939584e-05, 1.939584e-05, 
    1.939582e-05, 1.939581e-05, 1.93958e-05, 1.939579e-05, 1.939578e-05, 
    1.939576e-05, 1.939575e-05, 1.939572e-05, 1.939573e-05, 1.939572e-05, 
    1.939571e-05, 1.93957e-05, 1.93957e-05, 1.93957e-05, 1.939572e-05, 
    1.93957e-05, 1.939573e-05, 1.939572e-05, 1.939578e-05, 1.93958e-05, 
    1.939581e-05, 1.939582e-05, 1.939584e-05, 1.939583e-05, 1.939583e-05, 
    1.939582e-05, 1.939581e-05, 1.939581e-05, 1.939579e-05, 1.93958e-05, 
    1.939575e-05, 1.939577e-05, 1.939571e-05, 1.939573e-05, 1.939571e-05, 
    1.939572e-05, 1.93957e-05, 1.939572e-05, 1.939569e-05, 1.939569e-05, 
    1.939569e-05, 1.939568e-05, 1.939572e-05, 1.93957e-05, 1.939581e-05, 
    1.939581e-05, 1.939581e-05, 1.939583e-05, 1.939583e-05, 1.939584e-05, 
    1.939583e-05, 1.939582e-05, 1.939581e-05, 1.93958e-05, 1.93958e-05, 
    1.939578e-05, 1.939577e-05, 1.939574e-05, 1.939573e-05, 1.939571e-05, 
    1.939572e-05, 1.939572e-05, 1.939572e-05, 1.939573e-05, 1.939569e-05, 
    1.939571e-05, 1.939568e-05, 1.939568e-05, 1.93957e-05, 1.939568e-05, 
    1.939581e-05, 1.939582e-05, 1.939583e-05, 1.939582e-05, 1.939584e-05, 
    1.939583e-05, 1.939582e-05, 1.93958e-05, 1.939579e-05, 1.939579e-05, 
    1.939578e-05, 1.939577e-05, 1.939575e-05, 1.939573e-05, 1.939571e-05, 
    1.939571e-05, 1.939571e-05, 1.939571e-05, 1.939572e-05, 1.939571e-05, 
    1.939571e-05, 1.939571e-05, 1.939568e-05, 1.939569e-05, 1.939568e-05, 
    1.939569e-05, 1.939582e-05, 1.939581e-05, 1.939581e-05, 1.939581e-05, 
    1.939581e-05, 1.939579e-05, 1.939579e-05, 1.939576e-05, 1.939577e-05, 
    1.939575e-05, 1.939577e-05, 1.939576e-05, 1.939575e-05, 1.939577e-05, 
    1.939573e-05, 1.939575e-05, 1.939571e-05, 1.939573e-05, 1.939571e-05, 
    1.939571e-05, 1.93957e-05, 1.93957e-05, 1.939569e-05, 1.939567e-05, 
    1.939568e-05, 1.939566e-05, 1.93958e-05, 1.939579e-05, 1.939579e-05, 
    1.939578e-05, 1.939578e-05, 1.939576e-05, 1.939574e-05, 1.939575e-05, 
    1.939573e-05, 1.939573e-05, 1.939575e-05, 1.939574e-05, 1.939579e-05, 
    1.939578e-05, 1.939578e-05, 1.93958e-05, 1.939575e-05, 1.939577e-05, 
    1.939573e-05, 1.939574e-05, 1.93957e-05, 1.939572e-05, 1.939568e-05, 
    1.939566e-05, 1.939565e-05, 1.939563e-05, 1.939579e-05, 1.939579e-05, 
    1.939578e-05, 1.939577e-05, 1.939576e-05, 1.939574e-05, 1.939574e-05, 
    1.939573e-05, 1.939573e-05, 1.939572e-05, 1.939573e-05, 1.939572e-05, 
    1.939578e-05, 1.939575e-05, 1.93958e-05, 1.939578e-05, 1.939577e-05, 
    1.939577e-05, 1.939575e-05, 1.939575e-05, 1.939572e-05, 1.939573e-05, 
    1.939567e-05, 1.93957e-05, 1.939561e-05, 1.939563e-05, 1.939579e-05, 
    1.939579e-05, 1.939576e-05, 1.939577e-05, 1.939574e-05, 1.939573e-05, 
    1.939572e-05, 1.939571e-05, 1.939571e-05, 1.939571e-05, 1.939572e-05, 
    1.939571e-05, 1.939574e-05, 1.939573e-05, 1.939576e-05, 1.939575e-05, 
    1.939576e-05, 1.939576e-05, 1.939575e-05, 1.939573e-05, 1.939573e-05, 
    1.939573e-05, 1.939571e-05, 1.939574e-05, 1.939566e-05, 1.939571e-05, 
    1.939578e-05, 1.939577e-05, 1.939576e-05, 1.939577e-05, 1.939573e-05, 
    1.939574e-05, 1.939571e-05, 1.939572e-05, 1.93957e-05, 1.939571e-05, 
    1.939571e-05, 1.939572e-05, 1.939573e-05, 1.939574e-05, 1.939576e-05, 
    1.939577e-05, 1.939577e-05, 1.939575e-05, 1.939573e-05, 1.939571e-05, 
    1.939572e-05, 1.93957e-05, 1.939574e-05, 1.939572e-05, 1.939573e-05, 
    1.939571e-05, 1.939575e-05, 1.939572e-05, 1.939576e-05, 1.939575e-05, 
    1.939574e-05, 1.939572e-05, 1.939572e-05, 1.939571e-05, 1.939572e-05, 
    1.939573e-05, 1.939573e-05, 1.939575e-05, 1.939575e-05, 1.939576e-05, 
    1.939576e-05, 1.939576e-05, 1.939575e-05, 1.939573e-05, 1.939571e-05, 
    1.93957e-05, 1.939569e-05, 1.939567e-05, 1.939569e-05, 1.939566e-05, 
    1.939569e-05, 1.939564e-05, 1.939572e-05, 1.939569e-05, 1.939574e-05, 
    1.939574e-05, 1.939573e-05, 1.93957e-05, 1.939571e-05, 1.93957e-05, 
    1.939573e-05, 1.939575e-05, 1.939576e-05, 1.939577e-05, 1.939576e-05, 
    1.939576e-05, 1.939575e-05, 1.939575e-05, 1.939573e-05, 1.939574e-05, 
    1.939571e-05, 1.93957e-05, 1.939566e-05, 1.939564e-05, 1.939562e-05, 
    1.939561e-05, 1.939561e-05, 1.939561e-05 ;

 LITR2C_TO_SOIL1C =
  1.23344e-13, 1.236579e-13, 1.235969e-13, 1.238499e-13, 1.237097e-13, 
    1.238752e-13, 1.234077e-13, 1.236703e-13, 1.235027e-13, 1.233723e-13, 
    1.243401e-13, 1.238612e-13, 1.248371e-13, 1.245322e-13, 1.252974e-13, 
    1.247896e-13, 1.253997e-13, 1.252829e-13, 1.256346e-13, 1.255339e-13, 
    1.25983e-13, 1.256811e-13, 1.262157e-13, 1.25911e-13, 1.259587e-13, 
    1.256711e-13, 1.239578e-13, 1.242805e-13, 1.239386e-13, 1.239847e-13, 
    1.23964e-13, 1.237125e-13, 1.235856e-13, 1.2332e-13, 1.233683e-13, 
    1.235634e-13, 1.240054e-13, 1.238555e-13, 1.242333e-13, 1.242248e-13, 
    1.246447e-13, 1.244554e-13, 1.251603e-13, 1.249602e-13, 1.255381e-13, 
    1.253929e-13, 1.255313e-13, 1.254893e-13, 1.255318e-13, 1.253188e-13, 
    1.254101e-13, 1.252226e-13, 1.244908e-13, 1.247061e-13, 1.240636e-13, 
    1.236764e-13, 1.234192e-13, 1.232364e-13, 1.232623e-13, 1.233115e-13, 
    1.235645e-13, 1.238023e-13, 1.239833e-13, 1.241043e-13, 1.242235e-13, 
    1.245837e-13, 1.247744e-13, 1.252007e-13, 1.251239e-13, 1.25254e-13, 
    1.253784e-13, 1.25587e-13, 1.255527e-13, 1.256445e-13, 1.252507e-13, 
    1.255125e-13, 1.250801e-13, 1.251984e-13, 1.242555e-13, 1.238959e-13, 
    1.237426e-13, 1.236087e-13, 1.232821e-13, 1.235076e-13, 1.234188e-13, 
    1.236302e-13, 1.237645e-13, 1.236981e-13, 1.241076e-13, 1.239485e-13, 
    1.247857e-13, 1.244254e-13, 1.253639e-13, 1.251397e-13, 1.254176e-13, 
    1.252759e-13, 1.255187e-13, 1.253002e-13, 1.256787e-13, 1.257611e-13, 
    1.257048e-13, 1.25921e-13, 1.25288e-13, 1.255312e-13, 1.236962e-13, 
    1.237071e-13, 1.237575e-13, 1.235356e-13, 1.235221e-13, 1.233187e-13, 
    1.234997e-13, 1.235767e-13, 1.237723e-13, 1.238879e-13, 1.239977e-13, 
    1.24239e-13, 1.245082e-13, 1.248843e-13, 1.251542e-13, 1.25335e-13, 
    1.252242e-13, 1.25322e-13, 1.252126e-13, 1.251614e-13, 1.257302e-13, 
    1.254109e-13, 1.258899e-13, 1.258634e-13, 1.256467e-13, 1.258664e-13, 
    1.237147e-13, 1.236524e-13, 1.234358e-13, 1.236053e-13, 1.232965e-13, 
    1.234694e-13, 1.235687e-13, 1.239517e-13, 1.240359e-13, 1.241138e-13, 
    1.242677e-13, 1.244651e-13, 1.248109e-13, 1.251115e-13, 1.253857e-13, 
    1.253656e-13, 1.253727e-13, 1.254338e-13, 1.252822e-13, 1.254587e-13, 
    1.254883e-13, 1.254109e-13, 1.258599e-13, 1.257317e-13, 1.258629e-13, 
    1.257794e-13, 1.236726e-13, 1.237775e-13, 1.237208e-13, 1.238273e-13, 
    1.237523e-13, 1.240857e-13, 1.241856e-13, 1.246527e-13, 1.244612e-13, 
    1.24766e-13, 1.244922e-13, 1.245407e-13, 1.247758e-13, 1.24507e-13, 
    1.250949e-13, 1.246963e-13, 1.254362e-13, 1.250386e-13, 1.254611e-13, 
    1.253845e-13, 1.255114e-13, 1.256249e-13, 1.257677e-13, 1.260309e-13, 
    1.2597e-13, 1.2619e-13, 1.239337e-13, 1.240695e-13, 1.240576e-13, 
    1.241997e-13, 1.243048e-13, 1.245324e-13, 1.248969e-13, 1.247599e-13, 
    1.250115e-13, 1.250619e-13, 1.246798e-13, 1.249144e-13, 1.241604e-13, 
    1.242823e-13, 1.242098e-13, 1.239444e-13, 1.247914e-13, 1.24357e-13, 
    1.251586e-13, 1.249238e-13, 1.256087e-13, 1.252682e-13, 1.259365e-13, 
    1.262214e-13, 1.264896e-13, 1.268023e-13, 1.241437e-13, 1.240514e-13, 
    1.242167e-13, 1.244449e-13, 1.246568e-13, 1.249381e-13, 1.249669e-13, 
    1.250195e-13, 1.251559e-13, 1.252704e-13, 1.250361e-13, 1.252992e-13, 
    1.243104e-13, 1.248291e-13, 1.240165e-13, 1.242613e-13, 1.244315e-13, 
    1.24357e-13, 1.247443e-13, 1.248354e-13, 1.252056e-13, 1.250144e-13, 
    1.261511e-13, 1.256488e-13, 1.270404e-13, 1.266522e-13, 1.240192e-13, 
    1.241434e-13, 1.245752e-13, 1.243698e-13, 1.249569e-13, 1.251011e-13, 
    1.252184e-13, 1.253681e-13, 1.253843e-13, 1.25473e-13, 1.253277e-13, 
    1.254673e-13, 1.249387e-13, 1.251751e-13, 1.24526e-13, 1.24684e-13, 
    1.246114e-13, 1.245316e-13, 1.247778e-13, 1.250397e-13, 1.250455e-13, 
    1.251294e-13, 1.253655e-13, 1.249593e-13, 1.262156e-13, 1.254402e-13, 
    1.242788e-13, 1.245176e-13, 1.245519e-13, 1.244594e-13, 1.250867e-13, 
    1.248595e-13, 1.254709e-13, 1.253058e-13, 1.255762e-13, 1.254419e-13, 
    1.254221e-13, 1.252495e-13, 1.251419e-13, 1.248699e-13, 1.246485e-13, 
    1.244728e-13, 1.245137e-13, 1.247066e-13, 1.250558e-13, 1.253858e-13, 
    1.253135e-13, 1.255557e-13, 1.249143e-13, 1.251834e-13, 1.250794e-13, 
    1.253505e-13, 1.247562e-13, 1.25262e-13, 1.246268e-13, 1.246825e-13, 
    1.24855e-13, 1.252016e-13, 1.252784e-13, 1.253601e-13, 1.253097e-13, 
    1.250647e-13, 1.250246e-13, 1.248509e-13, 1.248028e-13, 1.246704e-13, 
    1.245607e-13, 1.246609e-13, 1.247661e-13, 1.250648e-13, 1.253337e-13, 
    1.256265e-13, 1.256981e-13, 1.260395e-13, 1.257615e-13, 1.262199e-13, 
    1.2583e-13, 1.265047e-13, 1.252915e-13, 1.258187e-13, 1.248629e-13, 
    1.249661e-13, 1.251525e-13, 1.255797e-13, 1.253492e-13, 1.256188e-13, 
    1.25023e-13, 1.247132e-13, 1.246331e-13, 1.244835e-13, 1.246366e-13, 
    1.246241e-13, 1.247705e-13, 1.247235e-13, 1.250747e-13, 1.248861e-13, 
    1.254216e-13, 1.256167e-13, 1.26167e-13, 1.265036e-13, 1.26846e-13, 
    1.26997e-13, 1.270429e-13, 1.270621e-13 ;

 LITR2C_vr =
  0.001107522, 0.001107521, 0.001107521, 0.001107521, 0.001107521, 
    0.001107521, 0.001107522, 0.001107521, 0.001107522, 0.001107522, 
    0.001107519, 0.001107521, 0.001107517, 0.001107518, 0.001107516, 
    0.001107517, 0.001107515, 0.001107516, 0.001107514, 0.001107515, 
    0.001107513, 0.001107514, 0.001107512, 0.001107513, 0.001107513, 
    0.001107514, 0.00110752, 0.001107519, 0.00110752, 0.00110752, 0.00110752, 
    0.001107521, 0.001107521, 0.001107522, 0.001107522, 0.001107522, 
    0.00110752, 0.001107521, 0.001107519, 0.001107519, 0.001107518, 
    0.001107518, 0.001107516, 0.001107517, 0.001107515, 0.001107515, 
    0.001107515, 0.001107515, 0.001107515, 0.001107515, 0.001107515, 
    0.001107516, 0.001107518, 0.001107518, 0.00110752, 0.001107521, 
    0.001107522, 0.001107523, 0.001107523, 0.001107522, 0.001107522, 
    0.001107521, 0.00110752, 0.00110752, 0.001107519, 0.001107518, 
    0.001107517, 0.001107516, 0.001107516, 0.001107516, 0.001107515, 
    0.001107514, 0.001107515, 0.001107514, 0.001107516, 0.001107515, 
    0.001107516, 0.001107516, 0.001107519, 0.00110752, 0.001107521, 
    0.001107521, 0.001107523, 0.001107522, 0.001107522, 0.001107521, 
    0.001107521, 0.001107521, 0.00110752, 0.00110752, 0.001107517, 
    0.001107519, 0.001107515, 0.001107516, 0.001107515, 0.001107516, 
    0.001107515, 0.001107516, 0.001107514, 0.001107514, 0.001107514, 
    0.001107513, 0.001107516, 0.001107515, 0.001107521, 0.001107521, 
    0.001107521, 0.001107522, 0.001107522, 0.001107522, 0.001107522, 
    0.001107521, 0.001107521, 0.00110752, 0.00110752, 0.001107519, 
    0.001107518, 0.001107517, 0.001107516, 0.001107515, 0.001107516, 
    0.001107515, 0.001107516, 0.001107516, 0.001107514, 0.001107515, 
    0.001107513, 0.001107514, 0.001107514, 0.001107514, 0.001107521, 
    0.001107521, 0.001107522, 0.001107521, 0.001107523, 0.001107522, 
    0.001107522, 0.00110752, 0.00110752, 0.00110752, 0.001107519, 
    0.001107518, 0.001107517, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107515, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107514, 0.001107514, 0.001107514, 0.001107514, 
    0.001107521, 0.001107521, 0.001107521, 0.001107521, 0.001107521, 
    0.00110752, 0.001107519, 0.001107518, 0.001107518, 0.001107517, 
    0.001107518, 0.001107518, 0.001107517, 0.001107518, 0.001107516, 
    0.001107518, 0.001107515, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107514, 0.001107514, 0.001107513, 0.001107513, 
    0.001107512, 0.00110752, 0.00110752, 0.00110752, 0.001107519, 
    0.001107519, 0.001107518, 0.001107517, 0.001107517, 0.001107516, 
    0.001107516, 0.001107518, 0.001107517, 0.001107519, 0.001107519, 
    0.001107519, 0.00110752, 0.001107517, 0.001107519, 0.001107516, 
    0.001107517, 0.001107514, 0.001107516, 0.001107513, 0.001107512, 
    0.001107511, 0.00110751, 0.001107519, 0.00110752, 0.001107519, 
    0.001107518, 0.001107518, 0.001107517, 0.001107517, 0.001107516, 
    0.001107516, 0.001107516, 0.001107516, 0.001107516, 0.001107519, 
    0.001107517, 0.00110752, 0.001107519, 0.001107519, 0.001107519, 
    0.001107517, 0.001107517, 0.001107516, 0.001107516, 0.001107513, 
    0.001107514, 0.001107509, 0.001107511, 0.00110752, 0.001107519, 
    0.001107518, 0.001107519, 0.001107517, 0.001107516, 0.001107516, 
    0.001107515, 0.001107515, 0.001107515, 0.001107515, 0.001107515, 
    0.001107517, 0.001107516, 0.001107518, 0.001107518, 0.001107518, 
    0.001107518, 0.001107517, 0.001107516, 0.001107516, 0.001107516, 
    0.001107515, 0.001107517, 0.001107512, 0.001107515, 0.001107519, 
    0.001107518, 0.001107518, 0.001107518, 0.001107516, 0.001107517, 
    0.001107515, 0.001107516, 0.001107515, 0.001107515, 0.001107515, 
    0.001107516, 0.001107516, 0.001107517, 0.001107518, 0.001107518, 
    0.001107518, 0.001107518, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107517, 0.001107516, 0.001107516, 0.001107515, 
    0.001107517, 0.001107516, 0.001107518, 0.001107518, 0.001107517, 
    0.001107516, 0.001107516, 0.001107515, 0.001107516, 0.001107516, 
    0.001107516, 0.001107517, 0.001107517, 0.001107518, 0.001107518, 
    0.001107518, 0.001107517, 0.001107516, 0.001107515, 0.001107514, 
    0.001107514, 0.001107513, 0.001107514, 0.001107512, 0.001107514, 
    0.001107511, 0.001107516, 0.001107514, 0.001107517, 0.001107517, 
    0.001107516, 0.001107514, 0.001107515, 0.001107514, 0.001107516, 
    0.001107518, 0.001107518, 0.001107518, 0.001107518, 0.001107518, 
    0.001107517, 0.001107518, 0.001107516, 0.001107517, 0.001107515, 
    0.001107514, 0.001107513, 0.001107511, 0.00110751, 0.00110751, 
    0.001107509, 0.001107509,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684241e-07, 2.684239e-07, 2.684239e-07, 2.684237e-07, 2.684238e-07, 
    2.684237e-07, 2.684241e-07, 2.684238e-07, 2.68424e-07, 2.684241e-07, 
    2.684233e-07, 2.684237e-07, 2.684229e-07, 2.684231e-07, 2.684225e-07, 
    2.684229e-07, 2.684224e-07, 2.684225e-07, 2.684222e-07, 2.684223e-07, 
    2.684219e-07, 2.684221e-07, 2.684217e-07, 2.68422e-07, 2.684219e-07, 
    2.684222e-07, 2.684236e-07, 2.684233e-07, 2.684236e-07, 2.684236e-07, 
    2.684236e-07, 2.684238e-07, 2.684239e-07, 2.684241e-07, 2.684241e-07, 
    2.684239e-07, 2.684235e-07, 2.684237e-07, 2.684234e-07, 2.684234e-07, 
    2.68423e-07, 2.684232e-07, 2.684226e-07, 2.684228e-07, 2.684223e-07, 
    2.684224e-07, 2.684223e-07, 2.684223e-07, 2.684223e-07, 2.684224e-07, 
    2.684224e-07, 2.684225e-07, 2.684232e-07, 2.68423e-07, 2.684235e-07, 
    2.684238e-07, 2.684241e-07, 2.684242e-07, 2.684242e-07, 2.684241e-07, 
    2.684239e-07, 2.684237e-07, 2.684236e-07, 2.684235e-07, 2.684234e-07, 
    2.684231e-07, 2.684229e-07, 2.684226e-07, 2.684226e-07, 2.684225e-07, 
    2.684224e-07, 2.684222e-07, 2.684222e-07, 2.684222e-07, 2.684225e-07, 
    2.684223e-07, 2.684226e-07, 2.684226e-07, 2.684233e-07, 2.684237e-07, 
    2.684238e-07, 2.684239e-07, 2.684242e-07, 2.68424e-07, 2.684241e-07, 
    2.684239e-07, 2.684238e-07, 2.684238e-07, 2.684235e-07, 2.684236e-07, 
    2.684229e-07, 2.684232e-07, 2.684224e-07, 2.684226e-07, 2.684224e-07, 
    2.684225e-07, 2.684223e-07, 2.684225e-07, 2.684222e-07, 2.684221e-07, 
    2.684221e-07, 2.684219e-07, 2.684225e-07, 2.684223e-07, 2.684238e-07, 
    2.684238e-07, 2.684238e-07, 2.684239e-07, 2.68424e-07, 2.684241e-07, 
    2.68424e-07, 2.684239e-07, 2.684237e-07, 2.684237e-07, 2.684236e-07, 
    2.684233e-07, 2.684231e-07, 2.684228e-07, 2.684226e-07, 2.684224e-07, 
    2.684225e-07, 2.684224e-07, 2.684225e-07, 2.684226e-07, 2.684221e-07, 
    2.684224e-07, 2.68422e-07, 2.68422e-07, 2.684222e-07, 2.68422e-07, 
    2.684238e-07, 2.684239e-07, 2.68424e-07, 2.684239e-07, 2.684241e-07, 
    2.68424e-07, 2.684239e-07, 2.684236e-07, 2.684235e-07, 2.684235e-07, 
    2.684233e-07, 2.684232e-07, 2.684229e-07, 2.684226e-07, 2.684224e-07, 
    2.684224e-07, 2.684224e-07, 2.684224e-07, 2.684225e-07, 2.684223e-07, 
    2.684223e-07, 2.684224e-07, 2.68422e-07, 2.684221e-07, 2.68422e-07, 
    2.684221e-07, 2.684238e-07, 2.684237e-07, 2.684238e-07, 2.684237e-07, 
    2.684238e-07, 2.684235e-07, 2.684234e-07, 2.68423e-07, 2.684232e-07, 
    2.684229e-07, 2.684232e-07, 2.684231e-07, 2.684229e-07, 2.684231e-07, 
    2.684226e-07, 2.68423e-07, 2.684224e-07, 2.684227e-07, 2.684223e-07, 
    2.684224e-07, 2.684223e-07, 2.684222e-07, 2.684221e-07, 2.684218e-07, 
    2.684219e-07, 2.684217e-07, 2.684236e-07, 2.684235e-07, 2.684235e-07, 
    2.684234e-07, 2.684233e-07, 2.684231e-07, 2.684228e-07, 2.684229e-07, 
    2.684227e-07, 2.684227e-07, 2.68423e-07, 2.684228e-07, 2.684234e-07, 
    2.684233e-07, 2.684234e-07, 2.684236e-07, 2.684229e-07, 2.684233e-07, 
    2.684226e-07, 2.684228e-07, 2.684222e-07, 2.684225e-07, 2.684219e-07, 
    2.684217e-07, 2.684214e-07, 2.684212e-07, 2.684234e-07, 2.684235e-07, 
    2.684234e-07, 2.684232e-07, 2.68423e-07, 2.684228e-07, 2.684228e-07, 
    2.684227e-07, 2.684226e-07, 2.684225e-07, 2.684227e-07, 2.684225e-07, 
    2.684233e-07, 2.684229e-07, 2.684235e-07, 2.684233e-07, 2.684232e-07, 
    2.684233e-07, 2.684229e-07, 2.684229e-07, 2.684226e-07, 2.684227e-07, 
    2.684217e-07, 2.684222e-07, 2.68421e-07, 2.684213e-07, 2.684235e-07, 
    2.684234e-07, 2.684231e-07, 2.684233e-07, 2.684228e-07, 2.684226e-07, 
    2.684225e-07, 2.684224e-07, 2.684224e-07, 2.684223e-07, 2.684224e-07, 
    2.684223e-07, 2.684228e-07, 2.684226e-07, 2.684231e-07, 2.68423e-07, 
    2.68423e-07, 2.684231e-07, 2.684229e-07, 2.684227e-07, 2.684227e-07, 
    2.684226e-07, 2.684224e-07, 2.684228e-07, 2.684217e-07, 2.684224e-07, 
    2.684233e-07, 2.684231e-07, 2.684231e-07, 2.684232e-07, 2.684226e-07, 
    2.684228e-07, 2.684223e-07, 2.684225e-07, 2.684222e-07, 2.684224e-07, 
    2.684224e-07, 2.684225e-07, 2.684226e-07, 2.684228e-07, 2.68423e-07, 
    2.684232e-07, 2.684231e-07, 2.68423e-07, 2.684227e-07, 2.684224e-07, 
    2.684224e-07, 2.684222e-07, 2.684228e-07, 2.684226e-07, 2.684226e-07, 
    2.684224e-07, 2.684229e-07, 2.684225e-07, 2.68423e-07, 2.68423e-07, 
    2.684228e-07, 2.684226e-07, 2.684225e-07, 2.684224e-07, 2.684225e-07, 
    2.684227e-07, 2.684227e-07, 2.684228e-07, 2.684229e-07, 2.68423e-07, 
    2.684231e-07, 2.68423e-07, 2.684229e-07, 2.684227e-07, 2.684224e-07, 
    2.684222e-07, 2.684221e-07, 2.684218e-07, 2.684221e-07, 2.684217e-07, 
    2.68422e-07, 2.684214e-07, 2.684225e-07, 2.68422e-07, 2.684228e-07, 
    2.684228e-07, 2.684226e-07, 2.684222e-07, 2.684224e-07, 2.684222e-07, 
    2.684227e-07, 2.68423e-07, 2.68423e-07, 2.684232e-07, 2.68423e-07, 
    2.68423e-07, 2.684229e-07, 2.68423e-07, 2.684227e-07, 2.684228e-07, 
    2.684224e-07, 2.684222e-07, 2.684217e-07, 2.684214e-07, 2.684212e-07, 
    2.68421e-07, 2.68421e-07, 2.68421e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -1.56858e-25, 1.764652e-25, -3.921449e-26, 9.313441e-26, 3.186177e-26, 
    1.446034e-25, -7.352717e-26, -7.352717e-27, 1.960724e-25, -1.56858e-25, 
    1.936215e-25, -9.803622e-26, -5.882173e-26, 1.936215e-25, -1.838179e-25, 
    6.127264e-26, -3.651849e-25, -1.274471e-25, -9.803622e-26, -3.676358e-26, 
    4.166539e-26, 6.862535e-26, -1.249962e-25, -2.205815e-25, -1.200944e-25, 
    -8.578169e-26, 1.274471e-25, -4.166539e-26, 1.225453e-26, 1.053889e-25, 
    -2.426396e-25, 1.715634e-25, 4.65672e-26, 1.02938e-25, 1.225453e-26, 
    -8.578169e-26, -3.357741e-25, -1.617598e-25, -3.921449e-26, 1.421525e-25, 
    -6.862535e-26, -1.29898e-25, -4.65672e-26, -2.695996e-26, 2.695996e-26, 
    8.578169e-26, -8.82326e-26, -1.249962e-25, 7.352717e-26, 1.642107e-25, 
    1.519561e-25, -2.794032e-25, -4.65672e-26, -1.151926e-25, 7.597807e-26, 
    -9.558531e-26, -1.225453e-25, -6.127264e-26, 1.715634e-25, -9.803622e-26, 
    -2.156797e-25, -6.617445e-26, -9.068351e-26, -1.715634e-25, 6.127264e-26, 
    -3.431268e-25, -2.009742e-25, 5.882173e-26, -3.676358e-26, 1.347998e-25, 
    -1.666616e-25, -1.54407e-25, 9.313441e-26, 1.642107e-25, -3.431268e-26, 
    5.882173e-26, -1.838179e-25, -7.842898e-26, -2.279342e-25, -7.352717e-26, 
    8.82326e-26, 9.558531e-26, 1.530638e-41, 2.573451e-25, 1.887197e-25, 
    1.740143e-25, -1.81367e-25, -1.02938e-25, 1.176435e-25, -3.284213e-25, 
    -1.347998e-25, -7.597807e-26, 1.81367e-25, -1.789161e-25, -1.470543e-26, 
    1.421525e-25, -9.558531e-26, 6.127264e-26, 1.078398e-25, 7.842898e-26, 
    -1.151926e-25, -1.200944e-25, 2.843051e-25, -3.921449e-26, 2.009742e-25, 
    1.56858e-25, 5.146902e-26, -2.156797e-25, -1.225453e-25, 9.558531e-26, 
    -3.186177e-26, 2.352869e-25, 6.617445e-26, -2.009742e-25, -2.524433e-25, 
    5.146902e-26, 5.882173e-26, 9.313441e-26, 1.078398e-25, -7.842898e-26, 
    5.146902e-26, -2.450906e-27, 6.862535e-26, 1.715634e-25, -1.053889e-25, 
    1.740143e-25, -1.151926e-25, -4.901811e-27, 4.65672e-26, -4.901811e-27, 
    1.02938e-25, -4.166539e-26, -2.695996e-26, 1.176435e-25, -1.617598e-25, 
    -1.715634e-26, 1.470543e-25, 6.372354e-26, 6.372354e-26, 2.622469e-25, 
    1.151926e-25, 2.450906e-27, -9.803622e-27, -1.127417e-25, 2.205815e-26, 
    2.181306e-25, 1.078398e-25, 2.475414e-25, -1.151926e-25, -1.960724e-26, 
    1.225453e-25, -1.470543e-25, -6.862535e-26, -2.450906e-27, 1.102908e-25, 
    1.004871e-25, 5.637083e-26, -1.495052e-25, 1.519561e-25, -9.068351e-26, 
    -3.431268e-26, 9.558531e-26, -2.230324e-25, -2.058761e-25, 1.911706e-25, 
    -8.82326e-26, -1.274471e-25, -1.347998e-25, -1.54407e-25, -4.65672e-26, 
    -2.450906e-25, -1.004871e-25, 2.720505e-25, 2.867559e-25, -7.352717e-27, 
    -4.65672e-26, -1.225453e-25, -1.764652e-25, -1.56858e-25, -2.132288e-25, 
    9.803622e-27, -7.352717e-27, -2.671487e-25, -1.053889e-25, -1.102908e-25, 
    1.519561e-25, 2.377378e-25, -4.901811e-26, -1.715634e-26, 1.530638e-41, 
    -4.41163e-26, 1.960724e-26, 1.960724e-25, -2.450906e-27, -2.205815e-26, 
    2.941087e-26, -8.578169e-26, -2.034252e-25, 1.740143e-25, -9.313441e-26, 
    -2.034252e-25, 2.450905e-26, 2.058761e-25, -5.391992e-26, -7.842898e-26, 
    1.691125e-25, -1.54407e-25, -1.078398e-25, -2.107779e-25, 2.941087e-26, 
    1.323489e-25, 7.107626e-26, -5.146902e-26, -1.421525e-25, -1.249962e-25, 
    2.499924e-25, -9.558531e-26, -3.186177e-26, 4.901811e-27, -1.127417e-25, 
    1.642107e-25, 1.470543e-26, -7.597807e-26, -6.372354e-26, 9.068351e-26, 
    -8.333079e-26, 2.499924e-25, -1.519561e-25, -1.29898e-25, -1.102908e-25, 
    7.352717e-27, -1.789161e-25, -1.960724e-26, -2.965596e-25, 4.901811e-27, 
    2.941087e-26, 1.617598e-25, 1.421525e-25, 4.901811e-26, -5.391992e-26, 
    -3.186177e-26, -6.862535e-26, 7.842898e-26, -1.225453e-26, -2.450906e-27, 
    -1.127417e-25, -1.789161e-25, 7.107626e-26, -4.901811e-26, -9.313441e-26, 
    -1.887197e-25, -4.41163e-26, -1.740143e-25, -1.838179e-25, -3.676358e-26, 
    -2.794032e-25, -5.146902e-26, 2.009742e-25, 4.166539e-26, 8.82326e-26, 
    -3.676358e-26, -1.960724e-25, -1.225453e-26, -1.102908e-25, 
    -1.519561e-25, 1.936215e-25, 2.352869e-25, 2.450905e-26, -5.146902e-26, 
    -6.617445e-26, 8.333079e-26, -3.798904e-25, 2.132288e-25, -2.450905e-26, 
    -6.127264e-26, 1.225453e-25, -9.803622e-26, 1.225453e-26, -1.54407e-25, 
    1.127417e-25, 1.789161e-25, -5.882173e-26, -5.637083e-26, -7.842898e-26, 
    8.82326e-26, -2.941087e-26, -1.715634e-26, -7.107626e-26, -1.691125e-25, 
    -1.078398e-25, -2.941087e-26, 7.352717e-26, -5.391992e-26, 1.887197e-25, 
    -1.593089e-25, 1.127417e-25, -8.578169e-26, -4.65672e-26, 3.186177e-26, 
    -8.82326e-26, -1.593089e-25, 2.695996e-26, 9.803622e-26, -1.078398e-25, 
    -9.803622e-27, 8.087988e-26, -2.794032e-25, -2.303851e-25, -1.102908e-25, 
    7.352717e-26, -2.990105e-25, -2.08327e-25, 1.053889e-25, -5.637083e-26, 
    -2.009742e-25, 1.372507e-25, 1.715634e-25, 1.838179e-25, 1.225453e-25, 
    -1.397016e-25, -3.921449e-26, 1.323489e-25, 6.372354e-26, -9.313441e-26, 
    1.764652e-25, 1.397016e-25, 1.225453e-26, -1.421525e-25, -3.921449e-26, 
    2.475414e-25, -5.637083e-26, -6.617445e-26, 3.431268e-26, 2.499924e-25, 
    -1.225453e-26, -4.730248e-25, -6.372354e-26, -1.004871e-25,
  2.676227e-32, 2.676224e-32, 2.676225e-32, 2.676223e-32, 2.676224e-32, 
    2.676223e-32, 2.676227e-32, 2.676224e-32, 2.676226e-32, 2.676227e-32, 
    2.676219e-32, 2.676223e-32, 2.676214e-32, 2.676217e-32, 2.676211e-32, 
    2.676215e-32, 2.67621e-32, 2.676211e-32, 2.676208e-32, 2.676209e-32, 
    2.676205e-32, 2.676207e-32, 2.676203e-32, 2.676205e-32, 2.676205e-32, 
    2.676207e-32, 2.676222e-32, 2.676219e-32, 2.676222e-32, 2.676222e-32, 
    2.676222e-32, 2.676224e-32, 2.676225e-32, 2.676227e-32, 2.676227e-32, 
    2.676225e-32, 2.676222e-32, 2.676223e-32, 2.67622e-32, 2.67622e-32, 
    2.676216e-32, 2.676218e-32, 2.676212e-32, 2.676214e-32, 2.676209e-32, 
    2.67621e-32, 2.676209e-32, 2.676209e-32, 2.676209e-32, 2.67621e-32, 
    2.67621e-32, 2.676211e-32, 2.676217e-32, 2.676216e-32, 2.676221e-32, 
    2.676224e-32, 2.676227e-32, 2.676228e-32, 2.676228e-32, 2.676228e-32, 
    2.676225e-32, 2.676223e-32, 2.676222e-32, 2.676221e-32, 2.67622e-32, 
    2.676217e-32, 2.676215e-32, 2.676212e-32, 2.676212e-32, 2.676211e-32, 
    2.67621e-32, 2.676208e-32, 2.676209e-32, 2.676208e-32, 2.676211e-32, 
    2.676209e-32, 2.676212e-32, 2.676212e-32, 2.676219e-32, 2.676223e-32, 
    2.676224e-32, 2.676225e-32, 2.676228e-32, 2.676226e-32, 2.676227e-32, 
    2.676225e-32, 2.676224e-32, 2.676224e-32, 2.676221e-32, 2.676222e-32, 
    2.676215e-32, 2.676218e-32, 2.67621e-32, 2.676212e-32, 2.67621e-32, 
    2.676211e-32, 2.676209e-32, 2.676211e-32, 2.676207e-32, 2.676207e-32, 
    2.676207e-32, 2.676205e-32, 2.676211e-32, 2.676209e-32, 2.676224e-32, 
    2.676224e-32, 2.676224e-32, 2.676226e-32, 2.676226e-32, 2.676227e-32, 
    2.676226e-32, 2.676225e-32, 2.676224e-32, 2.676223e-32, 2.676222e-32, 
    2.67622e-32, 2.676217e-32, 2.676214e-32, 2.676212e-32, 2.67621e-32, 
    2.676211e-32, 2.67621e-32, 2.676211e-32, 2.676212e-32, 2.676207e-32, 
    2.67621e-32, 2.676206e-32, 2.676206e-32, 2.676208e-32, 2.676206e-32, 
    2.676224e-32, 2.676225e-32, 2.676227e-32, 2.676225e-32, 2.676228e-32, 
    2.676226e-32, 2.676225e-32, 2.676222e-32, 2.676222e-32, 2.676221e-32, 
    2.676219e-32, 2.676218e-32, 2.676215e-32, 2.676212e-32, 2.67621e-32, 
    2.67621e-32, 2.67621e-32, 2.676209e-32, 2.676211e-32, 2.676209e-32, 
    2.676209e-32, 2.67621e-32, 2.676206e-32, 2.676207e-32, 2.676206e-32, 
    2.676207e-32, 2.676224e-32, 2.676224e-32, 2.676224e-32, 2.676223e-32, 
    2.676224e-32, 2.676221e-32, 2.67622e-32, 2.676216e-32, 2.676218e-32, 
    2.676215e-32, 2.676217e-32, 2.676217e-32, 2.676215e-32, 2.676217e-32, 
    2.676212e-32, 2.676216e-32, 2.676209e-32, 2.676213e-32, 2.676209e-32, 
    2.67621e-32, 2.676209e-32, 2.676208e-32, 2.676207e-32, 2.676204e-32, 
    2.676205e-32, 2.676203e-32, 2.676222e-32, 2.676221e-32, 2.676221e-32, 
    2.67622e-32, 2.676219e-32, 2.676217e-32, 2.676214e-32, 2.676215e-32, 
    2.676213e-32, 2.676213e-32, 2.676216e-32, 2.676214e-32, 2.67622e-32, 
    2.676219e-32, 2.67622e-32, 2.676222e-32, 2.676215e-32, 2.676219e-32, 
    2.676212e-32, 2.676214e-32, 2.676208e-32, 2.676211e-32, 2.676205e-32, 
    2.676203e-32, 2.676201e-32, 2.676198e-32, 2.67622e-32, 2.676221e-32, 
    2.67622e-32, 2.676218e-32, 2.676216e-32, 2.676214e-32, 2.676214e-32, 
    2.676213e-32, 2.676212e-32, 2.676211e-32, 2.676213e-32, 2.676211e-32, 
    2.676219e-32, 2.676215e-32, 2.676222e-32, 2.676219e-32, 2.676218e-32, 
    2.676219e-32, 2.676215e-32, 2.676214e-32, 2.676212e-32, 2.676213e-32, 
    2.676203e-32, 2.676208e-32, 2.676196e-32, 2.676199e-32, 2.676222e-32, 
    2.67622e-32, 2.676217e-32, 2.676219e-32, 2.676214e-32, 2.676212e-32, 
    2.676211e-32, 2.67621e-32, 2.67621e-32, 2.676209e-32, 2.67621e-32, 
    2.676209e-32, 2.676214e-32, 2.676212e-32, 2.676217e-32, 2.676216e-32, 
    2.676217e-32, 2.676217e-32, 2.676215e-32, 2.676213e-32, 2.676213e-32, 
    2.676212e-32, 2.67621e-32, 2.676214e-32, 2.676203e-32, 2.676209e-32, 
    2.676219e-32, 2.676217e-32, 2.676217e-32, 2.676218e-32, 2.676212e-32, 
    2.676214e-32, 2.676209e-32, 2.676211e-32, 2.676208e-32, 2.676209e-32, 
    2.676209e-32, 2.676211e-32, 2.676212e-32, 2.676214e-32, 2.676216e-32, 
    2.676218e-32, 2.676217e-32, 2.676216e-32, 2.676213e-32, 2.67621e-32, 
    2.676211e-32, 2.676209e-32, 2.676214e-32, 2.676212e-32, 2.676212e-32, 
    2.67621e-32, 2.676215e-32, 2.676211e-32, 2.676216e-32, 2.676216e-32, 
    2.676214e-32, 2.676212e-32, 2.676211e-32, 2.67621e-32, 2.676211e-32, 
    2.676213e-32, 2.676213e-32, 2.676214e-32, 2.676215e-32, 2.676216e-32, 
    2.676217e-32, 2.676216e-32, 2.676215e-32, 2.676213e-32, 2.67621e-32, 
    2.676208e-32, 2.676207e-32, 2.676204e-32, 2.676207e-32, 2.676203e-32, 
    2.676206e-32, 2.6762e-32, 2.676211e-32, 2.676206e-32, 2.676214e-32, 
    2.676214e-32, 2.676212e-32, 2.676208e-32, 2.67621e-32, 2.676208e-32, 
    2.676213e-32, 2.676216e-32, 2.676216e-32, 2.676218e-32, 2.676216e-32, 
    2.676217e-32, 2.676215e-32, 2.676216e-32, 2.676212e-32, 2.676214e-32, 
    2.676209e-32, 2.676208e-32, 2.676203e-32, 2.6762e-32, 2.676197e-32, 
    2.676196e-32, 2.676196e-32, 2.676196e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.413979e-15, 3.42267e-15, 3.420982e-15, 3.427984e-15, 3.424102e-15, 
    3.428685e-15, 3.415743e-15, 3.423013e-15, 3.418374e-15, 3.414764e-15, 
    3.44155e-15, 3.428297e-15, 3.455306e-15, 3.446869e-15, 3.468048e-15, 
    3.453992e-15, 3.47088e-15, 3.467646e-15, 3.477381e-15, 3.474594e-15, 
    3.487025e-15, 3.478668e-15, 3.493465e-15, 3.485032e-15, 3.48635e-15, 
    3.478391e-15, 3.430969e-15, 3.439901e-15, 3.430438e-15, 3.431713e-15, 
    3.431142e-15, 3.424181e-15, 3.420668e-15, 3.413317e-15, 3.414653e-15, 
    3.420053e-15, 3.432286e-15, 3.428138e-15, 3.438594e-15, 3.438359e-15, 
    3.449981e-15, 3.444743e-15, 3.464253e-15, 3.458714e-15, 3.47471e-15, 
    3.47069e-15, 3.474521e-15, 3.47336e-15, 3.474536e-15, 3.46864e-15, 
    3.471166e-15, 3.465976e-15, 3.445723e-15, 3.451681e-15, 3.433898e-15, 
    3.423181e-15, 3.416062e-15, 3.411004e-15, 3.411719e-15, 3.413082e-15, 
    3.420084e-15, 3.426665e-15, 3.431676e-15, 3.435025e-15, 3.438325e-15, 
    3.448294e-15, 3.453572e-15, 3.46537e-15, 3.463245e-15, 3.466847e-15, 
    3.47029e-15, 3.476064e-15, 3.475114e-15, 3.477656e-15, 3.466754e-15, 
    3.474e-15, 3.462034e-15, 3.465308e-15, 3.439211e-15, 3.429258e-15, 
    3.425014e-15, 3.421306e-15, 3.412269e-15, 3.41851e-15, 3.41605e-15, 
    3.421904e-15, 3.425619e-15, 3.423782e-15, 3.435117e-15, 3.430712e-15, 
    3.453884e-15, 3.443912e-15, 3.469889e-15, 3.463682e-15, 3.471376e-15, 
    3.467452e-15, 3.474174e-15, 3.468124e-15, 3.478603e-15, 3.480881e-15, 
    3.479324e-15, 3.485307e-15, 3.467788e-15, 3.47452e-15, 3.42373e-15, 
    3.42403e-15, 3.425427e-15, 3.419285e-15, 3.41891e-15, 3.41328e-15, 
    3.41829e-15, 3.420422e-15, 3.425836e-15, 3.429034e-15, 3.432074e-15, 
    3.438753e-15, 3.446204e-15, 3.456613e-15, 3.464084e-15, 3.469087e-15, 
    3.46602e-15, 3.468728e-15, 3.465701e-15, 3.464282e-15, 3.480027e-15, 
    3.471189e-15, 3.484447e-15, 3.483714e-15, 3.477716e-15, 3.483797e-15, 
    3.42424e-15, 3.422516e-15, 3.416523e-15, 3.421213e-15, 3.412667e-15, 
    3.417451e-15, 3.420199e-15, 3.430802e-15, 3.433132e-15, 3.435288e-15, 
    3.439549e-15, 3.445011e-15, 3.454583e-15, 3.462903e-15, 3.470491e-15, 
    3.469935e-15, 3.470131e-15, 3.471824e-15, 3.467628e-15, 3.472513e-15, 
    3.473331e-15, 3.47119e-15, 3.483616e-15, 3.480068e-15, 3.483699e-15, 
    3.481389e-15, 3.423077e-15, 3.425978e-15, 3.42441e-15, 3.427358e-15, 
    3.425281e-15, 3.43451e-15, 3.437275e-15, 3.450203e-15, 3.444903e-15, 
    3.453339e-15, 3.445761e-15, 3.447104e-15, 3.45361e-15, 3.446172e-15, 
    3.462442e-15, 3.451411e-15, 3.47189e-15, 3.460884e-15, 3.472579e-15, 
    3.470458e-15, 3.47397e-15, 3.477112e-15, 3.481065e-15, 3.488351e-15, 
    3.486665e-15, 3.492755e-15, 3.430303e-15, 3.434062e-15, 3.433733e-15, 
    3.437666e-15, 3.440573e-15, 3.446873e-15, 3.456963e-15, 3.453171e-15, 
    3.460133e-15, 3.461529e-15, 3.450953e-15, 3.457446e-15, 3.436578e-15, 
    3.439952e-15, 3.437945e-15, 3.430599e-15, 3.454042e-15, 3.442019e-15, 
    3.464207e-15, 3.457706e-15, 3.476664e-15, 3.46724e-15, 3.485736e-15, 
    3.493623e-15, 3.501047e-15, 3.509702e-15, 3.436115e-15, 3.433561e-15, 
    3.438134e-15, 3.444453e-15, 3.450317e-15, 3.458102e-15, 3.458899e-15, 
    3.460356e-15, 3.464131e-15, 3.467302e-15, 3.460815e-15, 3.468097e-15, 
    3.44073e-15, 3.455086e-15, 3.432594e-15, 3.439371e-15, 3.444082e-15, 
    3.442018e-15, 3.452738e-15, 3.455261e-15, 3.465507e-15, 3.460213e-15, 
    3.491676e-15, 3.477773e-15, 3.516291e-15, 3.505547e-15, 3.432669e-15, 
    3.436107e-15, 3.448058e-15, 3.442375e-15, 3.458623e-15, 3.462615e-15, 
    3.465862e-15, 3.470006e-15, 3.470454e-15, 3.472909e-15, 3.468886e-15, 
    3.472751e-15, 3.458119e-15, 3.464661e-15, 3.446695e-15, 3.451071e-15, 
    3.449059e-15, 3.44685e-15, 3.453666e-15, 3.460916e-15, 3.461074e-15, 
    3.463397e-15, 3.469933e-15, 3.458688e-15, 3.493462e-15, 3.472001e-15, 
    3.439854e-15, 3.446465e-15, 3.447412e-15, 3.444852e-15, 3.462215e-15, 
    3.455928e-15, 3.472849e-15, 3.468281e-15, 3.475766e-15, 3.472047e-15, 
    3.4715e-15, 3.466721e-15, 3.463743e-15, 3.456216e-15, 3.450086e-15, 
    3.445224e-15, 3.446355e-15, 3.451696e-15, 3.46136e-15, 3.470494e-15, 
    3.468493e-15, 3.475197e-15, 3.457446e-15, 3.464893e-15, 3.462014e-15, 
    3.469518e-15, 3.453069e-15, 3.467069e-15, 3.449485e-15, 3.451029e-15, 
    3.455803e-15, 3.465395e-15, 3.467521e-15, 3.469783e-15, 3.468388e-15, 
    3.461606e-15, 3.460496e-15, 3.455688e-15, 3.454359e-15, 3.450694e-15, 
    3.447656e-15, 3.450431e-15, 3.453342e-15, 3.46161e-15, 3.469051e-15, 
    3.477156e-15, 3.47914e-15, 3.488587e-15, 3.480893e-15, 3.493581e-15, 
    3.482789e-15, 3.501463e-15, 3.467884e-15, 3.482477e-15, 3.456022e-15, 
    3.458877e-15, 3.464036e-15, 3.475861e-15, 3.469483e-15, 3.476943e-15, 
    3.460453e-15, 3.451878e-15, 3.449662e-15, 3.445519e-15, 3.449757e-15, 
    3.449412e-15, 3.453465e-15, 3.452163e-15, 3.461885e-15, 3.456665e-15, 
    3.471485e-15, 3.476885e-15, 3.492116e-15, 3.501434e-15, 3.510912e-15, 
    3.51509e-15, 3.516362e-15, 3.516893e-15 ;

 LITR2N_vr =
  1.532729e-05, 1.532728e-05, 1.532728e-05, 1.532727e-05, 1.532728e-05, 
    1.532727e-05, 1.532729e-05, 1.532728e-05, 1.532729e-05, 1.532729e-05, 
    1.532725e-05, 1.532727e-05, 1.532722e-05, 1.532724e-05, 1.53272e-05, 
    1.532722e-05, 1.53272e-05, 1.53272e-05, 1.532718e-05, 1.532719e-05, 
    1.532717e-05, 1.532718e-05, 1.532716e-05, 1.532717e-05, 1.532717e-05, 
    1.532718e-05, 1.532726e-05, 1.532725e-05, 1.532726e-05, 1.532726e-05, 
    1.532726e-05, 1.532728e-05, 1.532728e-05, 1.53273e-05, 1.532729e-05, 
    1.532728e-05, 1.532726e-05, 1.532727e-05, 1.532725e-05, 1.532725e-05, 
    1.532723e-05, 1.532724e-05, 1.532721e-05, 1.532722e-05, 1.532719e-05, 
    1.53272e-05, 1.532719e-05, 1.532719e-05, 1.532719e-05, 1.53272e-05, 
    1.532719e-05, 1.53272e-05, 1.532724e-05, 1.532723e-05, 1.532726e-05, 
    1.532728e-05, 1.532729e-05, 1.53273e-05, 1.53273e-05, 1.53273e-05, 
    1.532728e-05, 1.532727e-05, 1.532726e-05, 1.532726e-05, 1.532725e-05, 
    1.532723e-05, 1.532722e-05, 1.53272e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.532719e-05, 1.532719e-05, 1.532718e-05, 1.53272e-05, 
    1.532719e-05, 1.532721e-05, 1.53272e-05, 1.532725e-05, 1.532727e-05, 
    1.532728e-05, 1.532728e-05, 1.53273e-05, 1.532729e-05, 1.532729e-05, 
    1.532728e-05, 1.532727e-05, 1.532728e-05, 1.532726e-05, 1.532726e-05, 
    1.532722e-05, 1.532724e-05, 1.53272e-05, 1.532721e-05, 1.532719e-05, 
    1.53272e-05, 1.532719e-05, 1.53272e-05, 1.532718e-05, 1.532718e-05, 
    1.532718e-05, 1.532717e-05, 1.53272e-05, 1.532719e-05, 1.532728e-05, 
    1.532728e-05, 1.532727e-05, 1.532728e-05, 1.532729e-05, 1.53273e-05, 
    1.532729e-05, 1.532728e-05, 1.532727e-05, 1.532727e-05, 1.532726e-05, 
    1.532725e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.53272e-05, 1.53272e-05, 1.532721e-05, 1.532718e-05, 
    1.532719e-05, 1.532717e-05, 1.532717e-05, 1.532718e-05, 1.532717e-05, 
    1.532728e-05, 1.532728e-05, 1.532729e-05, 1.532728e-05, 1.53273e-05, 
    1.532729e-05, 1.532728e-05, 1.532726e-05, 1.532726e-05, 1.532726e-05, 
    1.532725e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.53272e-05, 1.532719e-05, 1.53272e-05, 1.532719e-05, 
    1.532719e-05, 1.532719e-05, 1.532717e-05, 1.532718e-05, 1.532717e-05, 
    1.532718e-05, 1.532728e-05, 1.532727e-05, 1.532728e-05, 1.532727e-05, 
    1.532727e-05, 1.532726e-05, 1.532725e-05, 1.532723e-05, 1.532724e-05, 
    1.532722e-05, 1.532724e-05, 1.532724e-05, 1.532722e-05, 1.532724e-05, 
    1.532721e-05, 1.532723e-05, 1.532719e-05, 1.532721e-05, 1.532719e-05, 
    1.53272e-05, 1.532719e-05, 1.532718e-05, 1.532718e-05, 1.532716e-05, 
    1.532717e-05, 1.532716e-05, 1.532727e-05, 1.532726e-05, 1.532726e-05, 
    1.532725e-05, 1.532725e-05, 1.532724e-05, 1.532722e-05, 1.532723e-05, 
    1.532721e-05, 1.532721e-05, 1.532723e-05, 1.532722e-05, 1.532726e-05, 
    1.532725e-05, 1.532725e-05, 1.532726e-05, 1.532722e-05, 1.532724e-05, 
    1.532721e-05, 1.532722e-05, 1.532718e-05, 1.53272e-05, 1.532717e-05, 
    1.532716e-05, 1.532714e-05, 1.532713e-05, 1.532726e-05, 1.532726e-05, 
    1.532725e-05, 1.532724e-05, 1.532723e-05, 1.532722e-05, 1.532722e-05, 
    1.532721e-05, 1.532721e-05, 1.53272e-05, 1.532721e-05, 1.53272e-05, 
    1.532725e-05, 1.532722e-05, 1.532726e-05, 1.532725e-05, 1.532724e-05, 
    1.532724e-05, 1.532723e-05, 1.532722e-05, 1.53272e-05, 1.532721e-05, 
    1.532716e-05, 1.532718e-05, 1.532712e-05, 1.532713e-05, 1.532726e-05, 
    1.532726e-05, 1.532724e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 
    1.53272e-05, 1.53272e-05, 1.53272e-05, 1.532719e-05, 1.53272e-05, 
    1.532719e-05, 1.532722e-05, 1.532721e-05, 1.532724e-05, 1.532723e-05, 
    1.532723e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 1.532721e-05, 
    1.532721e-05, 1.53272e-05, 1.532722e-05, 1.532716e-05, 1.532719e-05, 
    1.532725e-05, 1.532724e-05, 1.532724e-05, 1.532724e-05, 1.532721e-05, 
    1.532722e-05, 1.532719e-05, 1.53272e-05, 1.532719e-05, 1.532719e-05, 
    1.532719e-05, 1.53272e-05, 1.532721e-05, 1.532722e-05, 1.532723e-05, 
    1.532724e-05, 1.532724e-05, 1.532723e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.532719e-05, 1.532722e-05, 1.53272e-05, 1.532721e-05, 
    1.53272e-05, 1.532723e-05, 1.53272e-05, 1.532723e-05, 1.532723e-05, 
    1.532722e-05, 1.53272e-05, 1.53272e-05, 1.53272e-05, 1.53272e-05, 
    1.532721e-05, 1.532721e-05, 1.532722e-05, 1.532722e-05, 1.532723e-05, 
    1.532724e-05, 1.532723e-05, 1.532722e-05, 1.532721e-05, 1.53272e-05, 
    1.532718e-05, 1.532718e-05, 1.532716e-05, 1.532718e-05, 1.532716e-05, 
    1.532717e-05, 1.532714e-05, 1.53272e-05, 1.532718e-05, 1.532722e-05, 
    1.532722e-05, 1.532721e-05, 1.532719e-05, 1.53272e-05, 1.532718e-05, 
    1.532721e-05, 1.532723e-05, 1.532723e-05, 1.532724e-05, 1.532723e-05, 
    1.532723e-05, 1.532722e-05, 1.532723e-05, 1.532721e-05, 1.532722e-05, 
    1.532719e-05, 1.532718e-05, 1.532716e-05, 1.532714e-05, 1.532712e-05, 
    1.532712e-05, 1.532712e-05, 1.532711e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.23344e-13, 1.236579e-13, 1.235969e-13, 1.238499e-13, 1.237097e-13, 
    1.238752e-13, 1.234077e-13, 1.236703e-13, 1.235027e-13, 1.233723e-13, 
    1.243401e-13, 1.238612e-13, 1.248371e-13, 1.245322e-13, 1.252974e-13, 
    1.247896e-13, 1.253997e-13, 1.252829e-13, 1.256346e-13, 1.255339e-13, 
    1.25983e-13, 1.256811e-13, 1.262157e-13, 1.25911e-13, 1.259587e-13, 
    1.256711e-13, 1.239578e-13, 1.242805e-13, 1.239386e-13, 1.239847e-13, 
    1.23964e-13, 1.237125e-13, 1.235856e-13, 1.2332e-13, 1.233683e-13, 
    1.235634e-13, 1.240054e-13, 1.238555e-13, 1.242333e-13, 1.242248e-13, 
    1.246447e-13, 1.244554e-13, 1.251603e-13, 1.249602e-13, 1.255381e-13, 
    1.253929e-13, 1.255313e-13, 1.254893e-13, 1.255318e-13, 1.253188e-13, 
    1.254101e-13, 1.252226e-13, 1.244908e-13, 1.247061e-13, 1.240636e-13, 
    1.236764e-13, 1.234192e-13, 1.232364e-13, 1.232623e-13, 1.233115e-13, 
    1.235645e-13, 1.238023e-13, 1.239833e-13, 1.241043e-13, 1.242235e-13, 
    1.245837e-13, 1.247744e-13, 1.252007e-13, 1.251239e-13, 1.25254e-13, 
    1.253784e-13, 1.25587e-13, 1.255527e-13, 1.256445e-13, 1.252507e-13, 
    1.255125e-13, 1.250801e-13, 1.251984e-13, 1.242555e-13, 1.238959e-13, 
    1.237426e-13, 1.236087e-13, 1.232821e-13, 1.235076e-13, 1.234188e-13, 
    1.236302e-13, 1.237645e-13, 1.236981e-13, 1.241076e-13, 1.239485e-13, 
    1.247857e-13, 1.244254e-13, 1.253639e-13, 1.251397e-13, 1.254176e-13, 
    1.252759e-13, 1.255187e-13, 1.253002e-13, 1.256787e-13, 1.257611e-13, 
    1.257048e-13, 1.25921e-13, 1.25288e-13, 1.255312e-13, 1.236962e-13, 
    1.237071e-13, 1.237575e-13, 1.235356e-13, 1.235221e-13, 1.233187e-13, 
    1.234997e-13, 1.235767e-13, 1.237723e-13, 1.238879e-13, 1.239977e-13, 
    1.24239e-13, 1.245082e-13, 1.248843e-13, 1.251542e-13, 1.25335e-13, 
    1.252242e-13, 1.25322e-13, 1.252126e-13, 1.251614e-13, 1.257302e-13, 
    1.254109e-13, 1.258899e-13, 1.258634e-13, 1.256467e-13, 1.258664e-13, 
    1.237147e-13, 1.236524e-13, 1.234358e-13, 1.236053e-13, 1.232965e-13, 
    1.234694e-13, 1.235687e-13, 1.239517e-13, 1.240359e-13, 1.241138e-13, 
    1.242677e-13, 1.244651e-13, 1.248109e-13, 1.251115e-13, 1.253857e-13, 
    1.253656e-13, 1.253727e-13, 1.254338e-13, 1.252822e-13, 1.254587e-13, 
    1.254883e-13, 1.254109e-13, 1.258599e-13, 1.257317e-13, 1.258629e-13, 
    1.257794e-13, 1.236726e-13, 1.237775e-13, 1.237208e-13, 1.238273e-13, 
    1.237523e-13, 1.240857e-13, 1.241856e-13, 1.246527e-13, 1.244612e-13, 
    1.24766e-13, 1.244922e-13, 1.245407e-13, 1.247758e-13, 1.24507e-13, 
    1.250949e-13, 1.246963e-13, 1.254362e-13, 1.250386e-13, 1.254611e-13, 
    1.253845e-13, 1.255114e-13, 1.256249e-13, 1.257677e-13, 1.260309e-13, 
    1.2597e-13, 1.2619e-13, 1.239337e-13, 1.240695e-13, 1.240576e-13, 
    1.241997e-13, 1.243048e-13, 1.245324e-13, 1.248969e-13, 1.247599e-13, 
    1.250115e-13, 1.250619e-13, 1.246798e-13, 1.249144e-13, 1.241604e-13, 
    1.242823e-13, 1.242098e-13, 1.239444e-13, 1.247914e-13, 1.24357e-13, 
    1.251586e-13, 1.249238e-13, 1.256087e-13, 1.252682e-13, 1.259365e-13, 
    1.262214e-13, 1.264896e-13, 1.268023e-13, 1.241437e-13, 1.240514e-13, 
    1.242167e-13, 1.244449e-13, 1.246568e-13, 1.249381e-13, 1.249669e-13, 
    1.250195e-13, 1.251559e-13, 1.252704e-13, 1.250361e-13, 1.252992e-13, 
    1.243104e-13, 1.248291e-13, 1.240165e-13, 1.242613e-13, 1.244315e-13, 
    1.24357e-13, 1.247443e-13, 1.248354e-13, 1.252056e-13, 1.250144e-13, 
    1.261511e-13, 1.256488e-13, 1.270404e-13, 1.266522e-13, 1.240192e-13, 
    1.241434e-13, 1.245752e-13, 1.243698e-13, 1.249569e-13, 1.251011e-13, 
    1.252184e-13, 1.253681e-13, 1.253843e-13, 1.25473e-13, 1.253277e-13, 
    1.254673e-13, 1.249387e-13, 1.251751e-13, 1.24526e-13, 1.24684e-13, 
    1.246114e-13, 1.245316e-13, 1.247778e-13, 1.250397e-13, 1.250455e-13, 
    1.251294e-13, 1.253655e-13, 1.249593e-13, 1.262156e-13, 1.254402e-13, 
    1.242788e-13, 1.245176e-13, 1.245519e-13, 1.244594e-13, 1.250867e-13, 
    1.248595e-13, 1.254709e-13, 1.253058e-13, 1.255762e-13, 1.254419e-13, 
    1.254221e-13, 1.252495e-13, 1.251419e-13, 1.248699e-13, 1.246485e-13, 
    1.244728e-13, 1.245137e-13, 1.247066e-13, 1.250558e-13, 1.253858e-13, 
    1.253135e-13, 1.255557e-13, 1.249143e-13, 1.251834e-13, 1.250794e-13, 
    1.253505e-13, 1.247562e-13, 1.25262e-13, 1.246268e-13, 1.246825e-13, 
    1.24855e-13, 1.252016e-13, 1.252784e-13, 1.253601e-13, 1.253097e-13, 
    1.250647e-13, 1.250246e-13, 1.248509e-13, 1.248028e-13, 1.246704e-13, 
    1.245607e-13, 1.246609e-13, 1.247661e-13, 1.250648e-13, 1.253337e-13, 
    1.256265e-13, 1.256981e-13, 1.260395e-13, 1.257615e-13, 1.262199e-13, 
    1.2583e-13, 1.265047e-13, 1.252915e-13, 1.258187e-13, 1.248629e-13, 
    1.249661e-13, 1.251525e-13, 1.255797e-13, 1.253492e-13, 1.256188e-13, 
    1.25023e-13, 1.247132e-13, 1.246331e-13, 1.244835e-13, 1.246366e-13, 
    1.246241e-13, 1.247705e-13, 1.247235e-13, 1.250747e-13, 1.248861e-13, 
    1.254216e-13, 1.256167e-13, 1.26167e-13, 1.265036e-13, 1.26846e-13, 
    1.26997e-13, 1.270429e-13, 1.270621e-13 ;

 LITR3C =
  9.697916e-06, 9.697906e-06, 9.697907e-06, 9.6979e-06, 9.697905e-06, 
    9.697899e-06, 9.697914e-06, 9.697906e-06, 9.697911e-06, 9.697915e-06, 
    9.697885e-06, 9.6979e-06, 9.69787e-06, 9.697879e-06, 9.697856e-06, 
    9.697871e-06, 9.697853e-06, 9.697857e-06, 9.697846e-06, 9.697848e-06, 
    9.697835e-06, 9.697844e-06, 9.697827e-06, 9.697837e-06, 9.697836e-06, 
    9.697845e-06, 9.697897e-06, 9.697887e-06, 9.697897e-06, 9.697896e-06, 
    9.697897e-06, 9.697905e-06, 9.697908e-06, 9.697917e-06, 9.697915e-06, 
    9.697909e-06, 9.697896e-06, 9.6979e-06, 9.697888e-06, 9.697888e-06, 
    9.697876e-06, 9.697882e-06, 9.69786e-06, 9.697867e-06, 9.697848e-06, 
    9.697853e-06, 9.697848e-06, 9.69785e-06, 9.697848e-06, 9.697856e-06, 
    9.697852e-06, 9.697858e-06, 9.69788e-06, 9.697874e-06, 9.697894e-06, 
    9.697906e-06, 9.697913e-06, 9.697919e-06, 9.697918e-06, 9.697917e-06, 
    9.697908e-06, 9.697901e-06, 9.697896e-06, 9.697892e-06, 9.697888e-06, 
    9.697877e-06, 9.697872e-06, 9.697859e-06, 9.697861e-06, 9.697857e-06, 
    9.697854e-06, 9.697847e-06, 9.697848e-06, 9.697846e-06, 9.697857e-06, 
    9.697849e-06, 9.697863e-06, 9.697859e-06, 9.697887e-06, 9.697898e-06, 
    9.697904e-06, 9.697907e-06, 9.697917e-06, 9.69791e-06, 9.697913e-06, 
    9.697907e-06, 9.697903e-06, 9.697905e-06, 9.697892e-06, 9.697897e-06, 
    9.697871e-06, 9.697883e-06, 9.697854e-06, 9.697861e-06, 9.697852e-06, 
    9.697857e-06, 9.697849e-06, 9.697856e-06, 9.697844e-06, 9.697842e-06, 
    9.697844e-06, 9.697837e-06, 9.697857e-06, 9.697848e-06, 9.697905e-06, 
    9.697905e-06, 9.697903e-06, 9.697909e-06, 9.69791e-06, 9.697917e-06, 
    9.697911e-06, 9.697908e-06, 9.697903e-06, 9.697899e-06, 9.697896e-06, 
    9.697888e-06, 9.69788e-06, 9.697868e-06, 9.69786e-06, 9.697855e-06, 
    9.697858e-06, 9.697855e-06, 9.697858e-06, 9.69786e-06, 9.697843e-06, 
    9.697852e-06, 9.697837e-06, 9.697838e-06, 9.697846e-06, 9.697838e-06, 
    9.697904e-06, 9.697907e-06, 9.697913e-06, 9.697907e-06, 9.697917e-06, 
    9.697912e-06, 9.697908e-06, 9.697897e-06, 9.697895e-06, 9.697892e-06, 
    9.697887e-06, 9.697881e-06, 9.697871e-06, 9.697862e-06, 9.697853e-06, 
    9.697854e-06, 9.697854e-06, 9.697852e-06, 9.697857e-06, 9.697851e-06, 
    9.69785e-06, 9.697852e-06, 9.697838e-06, 9.697843e-06, 9.697838e-06, 
    9.697841e-06, 9.697906e-06, 9.697902e-06, 9.697904e-06, 9.697901e-06, 
    9.697903e-06, 9.697893e-06, 9.69789e-06, 9.697876e-06, 9.697881e-06, 
    9.697872e-06, 9.69788e-06, 9.697879e-06, 9.697872e-06, 9.69788e-06, 
    9.697862e-06, 9.697874e-06, 9.697852e-06, 9.697864e-06, 9.697851e-06, 
    9.697853e-06, 9.697849e-06, 9.697846e-06, 9.697841e-06, 9.697834e-06, 
    9.697836e-06, 9.697828e-06, 9.697897e-06, 9.697894e-06, 9.697894e-06, 
    9.697889e-06, 9.697887e-06, 9.697879e-06, 9.697868e-06, 9.697872e-06, 
    9.697865e-06, 9.697863e-06, 9.697875e-06, 9.697867e-06, 9.69789e-06, 
    9.697887e-06, 9.697889e-06, 9.697897e-06, 9.697871e-06, 9.697885e-06, 
    9.69786e-06, 9.697867e-06, 9.697847e-06, 9.697857e-06, 9.697837e-06, 
    9.697827e-06, 9.697819e-06, 9.69781e-06, 9.697891e-06, 9.697894e-06, 
    9.697889e-06, 9.697882e-06, 9.697876e-06, 9.697867e-06, 9.697866e-06, 
    9.697865e-06, 9.69786e-06, 9.697857e-06, 9.697864e-06, 9.697856e-06, 
    9.697886e-06, 9.69787e-06, 9.697895e-06, 9.697887e-06, 9.697882e-06, 
    9.697885e-06, 9.697873e-06, 9.69787e-06, 9.697858e-06, 9.697865e-06, 
    9.69783e-06, 9.697845e-06, 9.697803e-06, 9.697815e-06, 9.697895e-06, 
    9.697891e-06, 9.697878e-06, 9.697884e-06, 9.697867e-06, 9.697862e-06, 
    9.697858e-06, 9.697854e-06, 9.697853e-06, 9.69785e-06, 9.697855e-06, 
    9.697851e-06, 9.697867e-06, 9.697859e-06, 9.697879e-06, 9.697875e-06, 
    9.697877e-06, 9.697879e-06, 9.697872e-06, 9.697864e-06, 9.697864e-06, 
    9.697861e-06, 9.697854e-06, 9.697867e-06, 9.697827e-06, 9.697851e-06, 
    9.697887e-06, 9.697879e-06, 9.697878e-06, 9.697881e-06, 9.697862e-06, 
    9.697869e-06, 9.69785e-06, 9.697856e-06, 9.697847e-06, 9.697851e-06, 
    9.697852e-06, 9.697857e-06, 9.69786e-06, 9.697869e-06, 9.697876e-06, 
    9.697881e-06, 9.69788e-06, 9.697874e-06, 9.697863e-06, 9.697853e-06, 
    9.697856e-06, 9.697848e-06, 9.697867e-06, 9.697859e-06, 9.697863e-06, 
    9.697854e-06, 9.697872e-06, 9.697857e-06, 9.697877e-06, 9.697875e-06, 
    9.697869e-06, 9.697858e-06, 9.697857e-06, 9.697854e-06, 9.697856e-06, 
    9.697863e-06, 9.697864e-06, 9.697869e-06, 9.697871e-06, 9.697875e-06, 
    9.697878e-06, 9.697876e-06, 9.697872e-06, 9.697863e-06, 9.697855e-06, 
    9.697846e-06, 9.697844e-06, 9.697833e-06, 9.697842e-06, 9.697827e-06, 
    9.697839e-06, 9.697819e-06, 9.697856e-06, 9.69784e-06, 9.697869e-06, 
    9.697866e-06, 9.69786e-06, 9.697847e-06, 9.697855e-06, 9.697846e-06, 
    9.697864e-06, 9.697874e-06, 9.697877e-06, 9.697881e-06, 9.697876e-06, 
    9.697877e-06, 9.697872e-06, 9.697874e-06, 9.697863e-06, 9.697868e-06, 
    9.697852e-06, 9.697847e-06, 9.697829e-06, 9.697819e-06, 9.697808e-06, 
    9.697804e-06, 9.697803e-06, 9.697802e-06 ;

 LITR3C_TO_SOIL2C =
  6.167196e-14, 6.182895e-14, 6.179845e-14, 6.192495e-14, 6.185481e-14, 
    6.19376e-14, 6.170383e-14, 6.183515e-14, 6.175134e-14, 6.168614e-14, 
    6.217002e-14, 6.19306e-14, 6.241851e-14, 6.22661e-14, 6.264869e-14, 
    6.239477e-14, 6.269984e-14, 6.264143e-14, 6.281729e-14, 6.276694e-14, 
    6.299149e-14, 6.284052e-14, 6.310782e-14, 6.295549e-14, 6.297931e-14, 
    6.283553e-14, 6.197886e-14, 6.214021e-14, 6.196928e-14, 6.199231e-14, 
    6.198199e-14, 6.185624e-14, 6.17928e-14, 6.165999e-14, 6.168412e-14, 
    6.178168e-14, 6.200266e-14, 6.192772e-14, 6.211662e-14, 6.211236e-14, 
    6.232231e-14, 6.222769e-14, 6.258012e-14, 6.248006e-14, 6.276904e-14, 
    6.269642e-14, 6.276562e-14, 6.274465e-14, 6.276589e-14, 6.265937e-14, 
    6.270502e-14, 6.261127e-14, 6.22454e-14, 6.235302e-14, 6.203178e-14, 
    6.183818e-14, 6.170958e-14, 6.16182e-14, 6.163113e-14, 6.165575e-14, 
    6.178224e-14, 6.190113e-14, 6.199164e-14, 6.205215e-14, 6.211175e-14, 
    6.229183e-14, 6.238717e-14, 6.260032e-14, 6.256193e-14, 6.262699e-14, 
    6.268919e-14, 6.279349e-14, 6.277634e-14, 6.282225e-14, 6.262531e-14, 
    6.275622e-14, 6.254004e-14, 6.25992e-14, 6.212775e-14, 6.194796e-14, 
    6.18713e-14, 6.180431e-14, 6.164106e-14, 6.175381e-14, 6.170937e-14, 
    6.181511e-14, 6.188223e-14, 6.184904e-14, 6.20538e-14, 6.197423e-14, 
    6.239283e-14, 6.221268e-14, 6.268194e-14, 6.256981e-14, 6.270881e-14, 
    6.263791e-14, 6.275935e-14, 6.265006e-14, 6.283936e-14, 6.288051e-14, 
    6.285238e-14, 6.296047e-14, 6.2644e-14, 6.27656e-14, 6.18481e-14, 
    6.185352e-14, 6.187875e-14, 6.17678e-14, 6.176102e-14, 6.165932e-14, 
    6.174983e-14, 6.178834e-14, 6.188614e-14, 6.194391e-14, 6.199883e-14, 
    6.211949e-14, 6.225408e-14, 6.244212e-14, 6.257708e-14, 6.266745e-14, 
    6.261206e-14, 6.266097e-14, 6.260629e-14, 6.258066e-14, 6.286508e-14, 
    6.270543e-14, 6.294493e-14, 6.29317e-14, 6.282334e-14, 6.293319e-14, 
    6.185732e-14, 6.182617e-14, 6.17179e-14, 6.180264e-14, 6.164824e-14, 
    6.173467e-14, 6.178432e-14, 6.197585e-14, 6.201794e-14, 6.20569e-14, 
    6.213386e-14, 6.223253e-14, 6.240544e-14, 6.255574e-14, 6.269282e-14, 
    6.268278e-14, 6.268631e-14, 6.27169e-14, 6.26411e-14, 6.272934e-14, 
    6.274413e-14, 6.270544e-14, 6.292992e-14, 6.286583e-14, 6.293141e-14, 
    6.288969e-14, 6.18363e-14, 6.188872e-14, 6.18604e-14, 6.191364e-14, 
    6.187612e-14, 6.204285e-14, 6.209279e-14, 6.232632e-14, 6.223058e-14, 
    6.238298e-14, 6.224608e-14, 6.227034e-14, 6.238787e-14, 6.22535e-14, 
    6.254742e-14, 6.234815e-14, 6.271809e-14, 6.251928e-14, 6.273053e-14, 
    6.269223e-14, 6.275566e-14, 6.281243e-14, 6.288384e-14, 6.301545e-14, 
    6.298499e-14, 6.3095e-14, 6.196684e-14, 6.203474e-14, 6.20288e-14, 
    6.209985e-14, 6.215236e-14, 6.226616e-14, 6.244844e-14, 6.237994e-14, 
    6.250571e-14, 6.253093e-14, 6.233986e-14, 6.245717e-14, 6.20802e-14, 
    6.214114e-14, 6.210488e-14, 6.197218e-14, 6.239567e-14, 6.217848e-14, 
    6.25793e-14, 6.246186e-14, 6.280433e-14, 6.263409e-14, 6.296821e-14, 
    6.311069e-14, 6.32448e-14, 6.340114e-14, 6.207183e-14, 6.20257e-14, 
    6.210831e-14, 6.222246e-14, 6.232838e-14, 6.246902e-14, 6.248342e-14, 
    6.250973e-14, 6.257792e-14, 6.263521e-14, 6.251802e-14, 6.264957e-14, 
    6.215519e-14, 6.241453e-14, 6.200823e-14, 6.213065e-14, 6.221575e-14, 
    6.217846e-14, 6.237211e-14, 6.24177e-14, 6.260278e-14, 6.250716e-14, 
    6.307551e-14, 6.282436e-14, 6.352017e-14, 6.332609e-14, 6.200957e-14, 
    6.207169e-14, 6.228758e-14, 6.21849e-14, 6.247842e-14, 6.255055e-14, 
    6.260919e-14, 6.268405e-14, 6.269215e-14, 6.273649e-14, 6.266383e-14, 
    6.273364e-14, 6.246932e-14, 6.258751e-14, 6.226296e-14, 6.234201e-14, 
    6.230566e-14, 6.226576e-14, 6.238888e-14, 6.251985e-14, 6.252271e-14, 
    6.256467e-14, 6.268274e-14, 6.247961e-14, 6.310778e-14, 6.27201e-14, 
    6.213937e-14, 6.225879e-14, 6.227592e-14, 6.222966e-14, 6.254332e-14, 
    6.242975e-14, 6.273542e-14, 6.265289e-14, 6.27881e-14, 6.272093e-14, 
    6.271104e-14, 6.262472e-14, 6.257093e-14, 6.243495e-14, 6.232422e-14, 
    6.223638e-14, 6.225681e-14, 6.235329e-14, 6.252788e-14, 6.269287e-14, 
    6.265673e-14, 6.277783e-14, 6.245716e-14, 6.259169e-14, 6.253969e-14, 
    6.267524e-14, 6.23781e-14, 6.2631e-14, 6.231336e-14, 6.234125e-14, 
    6.242749e-14, 6.260077e-14, 6.263916e-14, 6.268003e-14, 6.265482e-14, 
    6.253232e-14, 6.251226e-14, 6.242541e-14, 6.240139e-14, 6.233519e-14, 
    6.228032e-14, 6.233044e-14, 6.238303e-14, 6.253239e-14, 6.266681e-14, 
    6.281323e-14, 6.284905e-14, 6.301972e-14, 6.288072e-14, 6.310992e-14, 
    6.291497e-14, 6.325231e-14, 6.264573e-14, 6.290935e-14, 6.243144e-14, 
    6.248302e-14, 6.257621e-14, 6.278982e-14, 6.26746e-14, 6.280937e-14, 
    6.251148e-14, 6.235659e-14, 6.231655e-14, 6.224171e-14, 6.231826e-14, 
    6.231204e-14, 6.238525e-14, 6.236174e-14, 6.253735e-14, 6.244305e-14, 
    6.271078e-14, 6.280832e-14, 6.308346e-14, 6.325179e-14, 6.3423e-14, 
    6.349848e-14, 6.352145e-14, 6.353105e-14 ;

 LITR3C_vr =
  0.000553761, 0.0005537604, 0.0005537606, 0.0005537601, 0.0005537604, 
    0.0005537601, 0.0005537609, 0.0005537604, 0.0005537607, 0.000553761, 
    0.0005537593, 0.0005537601, 0.0005537584, 0.0005537589, 0.0005537576, 
    0.0005537585, 0.0005537574, 0.0005537576, 0.000553757, 0.0005537572, 
    0.0005537564, 0.0005537569, 0.000553756, 0.0005537565, 0.0005537564, 
    0.000553757, 0.0005537599, 0.0005537593, 0.00055376, 0.0005537599, 
    0.0005537599, 0.0005537603, 0.0005537606, 0.000553761, 0.000553761, 
    0.0005537606, 0.0005537599, 0.0005537601, 0.0005537595, 0.0005537595, 
    0.0005537588, 0.000553759, 0.0005537578, 0.0005537582, 0.0005537572, 
    0.0005537574, 0.0005537572, 0.0005537572, 0.0005537572, 0.0005537575, 
    0.0005537574, 0.0005537577, 0.000553759, 0.0005537586, 0.0005537597, 
    0.0005537604, 0.0005537609, 0.0005537612, 0.0005537611, 0.000553761, 
    0.0005537606, 0.0005537602, 0.0005537599, 0.0005537597, 0.0005537595, 
    0.0005537588, 0.0005537585, 0.0005537578, 0.0005537579, 0.0005537577, 
    0.0005537575, 0.0005537571, 0.0005537571, 0.000553757, 0.0005537577, 
    0.0005537572, 0.0005537579, 0.0005537578, 0.0005537594, 0.00055376, 
    0.0005537603, 0.0005537606, 0.0005537611, 0.0005537607, 0.0005537609, 
    0.0005537605, 0.0005537603, 0.0005537604, 0.0005537597, 0.0005537599, 
    0.0005537585, 0.0005537591, 0.0005537575, 0.0005537579, 0.0005537574, 
    0.0005537577, 0.0005537572, 0.0005537576, 0.000553757, 0.0005537568, 
    0.0005537569, 0.0005537565, 0.0005537576, 0.0005537572, 0.0005537604, 
    0.0005537604, 0.0005537603, 0.0005537607, 0.0005537607, 0.000553761, 
    0.0005537607, 0.0005537606, 0.0005537603, 0.00055376, 0.0005537599, 
    0.0005537595, 0.000553759, 0.0005537583, 0.0005537578, 0.0005537575, 
    0.0005537577, 0.0005537575, 0.0005537577, 0.0005537578, 0.0005537568, 
    0.0005537574, 0.0005537565, 0.0005537566, 0.000553757, 0.0005537566, 
    0.0005537603, 0.0005537604, 0.0005537609, 0.0005537606, 0.0005537611, 
    0.0005537608, 0.0005537606, 0.0005537599, 0.0005537598, 0.0005537596, 
    0.0005537594, 0.000553759, 0.0005537585, 0.0005537579, 0.0005537574, 
    0.0005537575, 0.0005537575, 0.0005537574, 0.0005537576, 0.0005537573, 
    0.0005537572, 0.0005537574, 0.0005537566, 0.0005537568, 0.0005537566, 
    0.0005537567, 0.0005537604, 0.0005537603, 0.0005537603, 0.0005537602, 
    0.0005537603, 0.0005537597, 0.0005537595, 0.0005537587, 0.000553759, 
    0.0005537585, 0.000553759, 0.0005537589, 0.0005537585, 0.000553759, 
    0.0005537579, 0.0005537586, 0.0005537574, 0.0005537581, 0.0005537573, 
    0.0005537574, 0.0005537572, 0.000553757, 0.0005537568, 0.0005537563, 
    0.0005537564, 0.000553756, 0.00055376, 0.0005537597, 0.0005537597, 
    0.0005537595, 0.0005537593, 0.0005537589, 0.0005537583, 0.0005537585, 
    0.0005537581, 0.000553758, 0.0005537586, 0.0005537582, 0.0005537596, 
    0.0005537593, 0.0005537595, 0.00055376, 0.0005537585, 0.0005537592, 
    0.0005537578, 0.0005537582, 0.0005537571, 0.0005537577, 0.0005537565, 
    0.000553756, 0.0005537555, 0.000553755, 0.0005537596, 0.0005537597, 
    0.0005537595, 0.0005537591, 0.0005537587, 0.0005537582, 0.0005537582, 
    0.0005537581, 0.0005537578, 0.0005537577, 0.0005537581, 0.0005537576, 
    0.0005537593, 0.0005537584, 0.0005537598, 0.0005537594, 0.0005537591, 
    0.0005537592, 0.0005537586, 0.0005537584, 0.0005537578, 0.0005537581, 
    0.0005537561, 0.000553757, 0.0005537546, 0.0005537552, 0.0005537598, 
    0.0005537596, 0.0005537589, 0.0005537592, 0.0005537582, 0.0005537579, 
    0.0005537577, 0.0005537575, 0.0005537574, 0.0005537573, 0.0005537575, 
    0.0005537573, 0.0005537582, 0.0005537578, 0.0005537589, 0.0005537586, 
    0.0005537588, 0.0005537589, 0.0005537585, 0.0005537581, 0.0005537581, 
    0.0005537579, 0.0005537575, 0.0005537582, 0.000553756, 0.0005537574, 
    0.0005537593, 0.0005537589, 0.0005537589, 0.000553759, 0.0005537579, 
    0.0005537583, 0.0005537573, 0.0005537576, 0.0005537571, 0.0005537574, 
    0.0005537574, 0.0005537577, 0.0005537579, 0.0005537583, 0.0005537587, 
    0.000553759, 0.0005537589, 0.0005537586, 0.000553758, 0.0005537574, 
    0.0005537575, 0.0005537571, 0.0005537582, 0.0005537578, 0.0005537579, 
    0.0005537575, 0.0005537585, 0.0005537577, 0.0005537588, 0.0005537586, 
    0.0005537583, 0.0005537578, 0.0005537577, 0.0005537575, 0.0005537576, 
    0.000553758, 0.0005537581, 0.0005537583, 0.0005537585, 0.0005537587, 
    0.0005537589, 0.0005537587, 0.0005537585, 0.000553758, 0.0005537575, 
    0.000553757, 0.0005537569, 0.0005537563, 0.0005537568, 0.000553756, 
    0.0005537567, 0.0005537555, 0.0005537576, 0.0005537567, 0.0005537583, 
    0.0005537582, 0.0005537578, 0.0005537571, 0.0005537575, 0.000553757, 
    0.0005537581, 0.0005537586, 0.0005537588, 0.000553759, 0.0005537588, 
    0.0005537588, 0.0005537585, 0.0005537586, 0.000553758, 0.0005537583, 
    0.0005537574, 0.000553757, 0.0005537561, 0.0005537555, 0.0005537549, 
    0.0005537546, 0.0005537546, 0.0005537545,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342121e-07, 1.342119e-07, 1.342119e-07, 1.342118e-07, 1.342119e-07, 
    1.342118e-07, 1.34212e-07, 1.342119e-07, 1.34212e-07, 1.34212e-07, 
    1.342116e-07, 1.342118e-07, 1.342114e-07, 1.342115e-07, 1.342112e-07, 
    1.342114e-07, 1.342112e-07, 1.342112e-07, 1.342111e-07, 1.342111e-07, 
    1.342109e-07, 1.342111e-07, 1.342108e-07, 1.34211e-07, 1.342109e-07, 
    1.342111e-07, 1.342118e-07, 1.342117e-07, 1.342118e-07, 1.342118e-07, 
    1.342118e-07, 1.342119e-07, 1.342119e-07, 1.342121e-07, 1.34212e-07, 
    1.34212e-07, 1.342118e-07, 1.342118e-07, 1.342117e-07, 1.342117e-07, 
    1.342115e-07, 1.342116e-07, 1.342113e-07, 1.342114e-07, 1.342111e-07, 
    1.342112e-07, 1.342111e-07, 1.342111e-07, 1.342111e-07, 1.342112e-07, 
    1.342112e-07, 1.342113e-07, 1.342116e-07, 1.342115e-07, 1.342117e-07, 
    1.342119e-07, 1.34212e-07, 1.342121e-07, 1.342121e-07, 1.342121e-07, 
    1.34212e-07, 1.342119e-07, 1.342118e-07, 1.342117e-07, 1.342117e-07, 
    1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342111e-07, 1.342111e-07, 1.342111e-07, 1.342112e-07, 
    1.342111e-07, 1.342113e-07, 1.342113e-07, 1.342117e-07, 1.342118e-07, 
    1.342119e-07, 1.342119e-07, 1.342121e-07, 1.34212e-07, 1.34212e-07, 
    1.342119e-07, 1.342119e-07, 1.342119e-07, 1.342117e-07, 1.342118e-07, 
    1.342114e-07, 1.342116e-07, 1.342112e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342111e-07, 1.342112e-07, 1.342111e-07, 1.34211e-07, 
    1.34211e-07, 1.34211e-07, 1.342112e-07, 1.342111e-07, 1.342119e-07, 
    1.342119e-07, 1.342119e-07, 1.34212e-07, 1.34212e-07, 1.342121e-07, 
    1.34212e-07, 1.34212e-07, 1.342119e-07, 1.342118e-07, 1.342118e-07, 
    1.342117e-07, 1.342116e-07, 1.342114e-07, 1.342113e-07, 1.342112e-07, 
    1.342113e-07, 1.342112e-07, 1.342113e-07, 1.342113e-07, 1.34211e-07, 
    1.342112e-07, 1.34211e-07, 1.34211e-07, 1.342111e-07, 1.34211e-07, 
    1.342119e-07, 1.342119e-07, 1.34212e-07, 1.342119e-07, 1.342121e-07, 
    1.34212e-07, 1.34212e-07, 1.342118e-07, 1.342118e-07, 1.342117e-07, 
    1.342117e-07, 1.342116e-07, 1.342114e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342112e-07, 1.342112e-07, 1.342112e-07, 1.342112e-07, 
    1.342111e-07, 1.342112e-07, 1.34211e-07, 1.34211e-07, 1.34211e-07, 
    1.34211e-07, 1.342119e-07, 1.342119e-07, 1.342119e-07, 1.342118e-07, 
    1.342119e-07, 1.342117e-07, 1.342117e-07, 1.342115e-07, 1.342116e-07, 
    1.342114e-07, 1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342116e-07, 
    1.342113e-07, 1.342115e-07, 1.342112e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342111e-07, 1.342111e-07, 1.34211e-07, 1.342109e-07, 
    1.342109e-07, 1.342109e-07, 1.342118e-07, 1.342117e-07, 1.342117e-07, 
    1.342117e-07, 1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342114e-07, 
    1.342113e-07, 1.342113e-07, 1.342115e-07, 1.342114e-07, 1.342117e-07, 
    1.342117e-07, 1.342117e-07, 1.342118e-07, 1.342114e-07, 1.342116e-07, 
    1.342113e-07, 1.342114e-07, 1.342111e-07, 1.342112e-07, 1.342109e-07, 
    1.342108e-07, 1.342107e-07, 1.342106e-07, 1.342117e-07, 1.342118e-07, 
    1.342117e-07, 1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342114e-07, 
    1.342113e-07, 1.342113e-07, 1.342112e-07, 1.342113e-07, 1.342112e-07, 
    1.342116e-07, 1.342114e-07, 1.342118e-07, 1.342117e-07, 1.342116e-07, 
    1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 
    1.342109e-07, 1.342111e-07, 1.342105e-07, 1.342107e-07, 1.342118e-07, 
    1.342117e-07, 1.342115e-07, 1.342116e-07, 1.342114e-07, 1.342113e-07, 
    1.342113e-07, 1.342112e-07, 1.342112e-07, 1.342111e-07, 1.342112e-07, 
    1.342111e-07, 1.342114e-07, 1.342113e-07, 1.342115e-07, 1.342115e-07, 
    1.342115e-07, 1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 
    1.342113e-07, 1.342112e-07, 1.342114e-07, 1.342108e-07, 1.342112e-07, 
    1.342117e-07, 1.342116e-07, 1.342115e-07, 1.342116e-07, 1.342113e-07, 
    1.342114e-07, 1.342111e-07, 1.342112e-07, 1.342111e-07, 1.342112e-07, 
    1.342112e-07, 1.342112e-07, 1.342113e-07, 1.342114e-07, 1.342115e-07, 
    1.342116e-07, 1.342116e-07, 1.342115e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342111e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 
    1.342112e-07, 1.342115e-07, 1.342112e-07, 1.342115e-07, 1.342115e-07, 
    1.342114e-07, 1.342113e-07, 1.342112e-07, 1.342112e-07, 1.342112e-07, 
    1.342113e-07, 1.342113e-07, 1.342114e-07, 1.342114e-07, 1.342115e-07, 
    1.342115e-07, 1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342112e-07, 
    1.342111e-07, 1.342111e-07, 1.342109e-07, 1.34211e-07, 1.342108e-07, 
    1.34211e-07, 1.342107e-07, 1.342112e-07, 1.34211e-07, 1.342114e-07, 
    1.342114e-07, 1.342113e-07, 1.342111e-07, 1.342112e-07, 1.342111e-07, 
    1.342113e-07, 1.342115e-07, 1.342115e-07, 1.342116e-07, 1.342115e-07, 
    1.342115e-07, 1.342114e-07, 1.342115e-07, 1.342113e-07, 1.342114e-07, 
    1.342112e-07, 1.342111e-07, 1.342109e-07, 1.342107e-07, 1.342106e-07, 
    1.342105e-07, 1.342105e-07, 1.342105e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  -1.017126e-25, 4.534175e-26, -7.352717e-27, -2.08327e-26, 5.146902e-26, 
    -1.960724e-26, -3.921449e-26, 1.409271e-25, -4.65672e-26, -9.068351e-26, 
    1.139671e-25, -7.352717e-26, -3.676358e-27, 1.960724e-26, -6.127264e-26, 
    2.08327e-26, -4.534175e-26, 3.431268e-26, 9.803622e-27, -3.186177e-26, 
    3.798904e-26, -6.4949e-26, -3.676358e-26, -4.043994e-26, 1.372507e-25, 
    2.205815e-26, 1.017126e-25, -1.004871e-25, -4.166539e-26, -3.308722e-26, 
    -9.803622e-27, -1.838179e-26, -2.818541e-26, 3.676358e-26, 1.102908e-26, 
    6.98508e-26, -5.637083e-26, 2.695996e-26, 2.573451e-26, 5.637083e-26, 
    -4.043994e-26, -8.087988e-26, 4.41163e-26, 9.313441e-26, 6.617445e-26, 
    8.82326e-26, -5.269447e-26, 7.965443e-26, 7.352717e-27, -6.127264e-26, 
    4.901811e-27, 5.269447e-26, -5.146902e-26, 4.65672e-26, 1.311234e-25, 
    5.146902e-26, -2.941087e-26, 7.352717e-27, 3.798904e-26, 1.090653e-25, 
    -5.514538e-26, -4.41163e-26, 5.637083e-26, -4.901811e-27, -4.901811e-26, 
    -2.205815e-26, -1.053889e-25, 6.73999e-26, -1.727888e-25, -7.352717e-27, 
    3.308722e-26, -4.166539e-26, 1.81367e-25, -1.090653e-25, -6.127264e-27, 
    4.41163e-26, -2.941087e-26, 4.534175e-26, 1.470543e-26, 2.450905e-26, 
    3.553813e-26, -6.617445e-26, 6.127264e-26, -6.4949e-26, 2.450905e-26, 
    -9.803622e-26, -1.593089e-26, 4.41163e-26, -1.347998e-26, -6.862535e-26, 
    1.56858e-25, -2.818541e-26, 7.965443e-26, -1.470543e-26, -8.578169e-27, 
    -3.308722e-26, 7.652491e-42, 4.901811e-27, 5.146902e-26, -5.759628e-26, 
    -1.531816e-25, 6.617445e-26, -2.941087e-26, 1.960724e-25, -9.803622e-27, 
    8.210533e-26, -4.043994e-26, 7.720352e-26, 5.269447e-26, -8.82326e-26, 
    -8.578169e-26, -6.127264e-26, -1.960724e-26, -4.41163e-26, -1.715634e-26, 
    -1.041635e-25, 4.901811e-27, 3.063632e-26, 6.73999e-26, -3.553813e-26, 
    -3.676358e-27, 2.695996e-26, 4.289085e-26, -4.901811e-27, -2.695996e-26, 
    4.901811e-27, 4.166539e-26, 1.409271e-25, 2.205815e-26, 3.921449e-26, 
    1.593089e-26, 1.556325e-25, 4.289085e-26, 7.107626e-26, -7.352717e-27, 
    4.043994e-26, -7.230172e-26, -3.186177e-26, 4.043994e-26, -1.200944e-25, 
    -4.901811e-27, -6.4949e-26, 8.087988e-26, 9.803622e-27, 2.450906e-27, 
    1.715634e-26, 4.65672e-26, -8.578169e-26, 4.289085e-26, 8.455624e-26, 
    4.534175e-26, -7.352717e-27, -5.146902e-26, -1.347998e-26, 6.372354e-26, 
    8.087988e-26, 1.960724e-26, -1.02938e-25, -6.127264e-26, 7.352717e-27, 
    -6.98508e-26, -7.597807e-26, 8.945805e-26, -5.882173e-26, 9.313441e-26, 
    -7.597807e-26, 7.652491e-42, 7.720352e-26, 1.470543e-25, 4.901811e-26, 
    6.127264e-27, -6.249809e-26, -9.926167e-26, 4.41163e-26, 1.176435e-25, 
    -2.450905e-26, 4.534175e-26, 1.593089e-26, 1.115162e-25, -8.087988e-26, 
    -3.186177e-26, -6.004719e-26, -4.901811e-27, 2.303851e-25, 2.08327e-26, 
    7.842898e-26, -7.475262e-26, 1.838179e-26, -3.431268e-26, -5.637083e-26, 
    0, 1.470543e-26, 6.862535e-26, 1.262216e-25, -5.269447e-26, 5.391992e-26, 
    -3.431268e-26, 7.352717e-26, 2.156797e-25, -5.024356e-26, 3.308722e-26, 
    1.225453e-27, 4.166539e-26, 8.210533e-26, 2.205815e-26, -1.078398e-25, 
    5.146902e-26, -4.043994e-26, -2.450906e-27, -4.043994e-26, -8.578169e-26, 
    8.210533e-26, 1.225453e-26, -2.818541e-26, -6.73999e-26, -7.965443e-26, 
    1.053889e-25, -1.347998e-26, 7.842898e-26, -1.642107e-25, -1.102908e-26, 
    -6.004719e-26, -2.450906e-27, -2.941087e-26, -3.676358e-27, 
    -4.779266e-26, 1.213198e-25, -5.637083e-26, -1.311234e-25, 9.558531e-26, 
    1.237707e-25, 3.431268e-26, -3.063632e-26, 8.333079e-26, 5.637083e-26, 
    1.593089e-26, 1.225453e-27, 5.514538e-26, 1.237707e-25, 1.593089e-26, 
    3.676358e-26, 9.803622e-26, 4.534175e-26, -5.391992e-26, -1.838179e-26, 
    -4.043994e-26, 1.225453e-26, -8.578169e-27, -4.289085e-26, -2.818541e-26, 
    2.941087e-26, -5.637083e-26, -2.205815e-26, 1.225453e-25, -2.695996e-26, 
    -9.803622e-27, 7.230172e-26, -4.043994e-26, 8.945805e-26, 1.960724e-26, 
    -6.73999e-26, -3.431268e-26, -1.102908e-26, 8.700715e-26, 3.186177e-26, 
    2.205815e-26, 5.391992e-26, 3.308722e-26, 2.573451e-26, 1.384762e-25, 
    1.16418e-25, -8.455624e-26, -1.838179e-26, -6.73999e-26, -5.882173e-26, 
    4.41163e-26, -4.65672e-26, -6.98508e-26, -5.514538e-26, -3.676358e-26, 
    2.450905e-26, -5.024356e-26, -7.352717e-26, -1.470543e-26, -2.818541e-26, 
    -6.372354e-26, -1.188689e-25, -1.335744e-25, 1.347998e-26, -9.313441e-26, 
    -2.450906e-27, -4.166539e-26, -3.798904e-26, -4.901811e-27, 1.960724e-26, 
    2.450906e-27, 2.818541e-26, 9.803622e-26, 4.043994e-26, 1.838179e-26, 
    -2.941087e-26, -6.372354e-26, -4.41163e-26, -1.715634e-26, 5.269447e-26, 
    -1.102908e-26, -3.676358e-26, 1.960724e-26, 4.65672e-26, 9.803622e-27, 
    -6.127264e-27, 1.642107e-25, -7.965443e-26, -7.352717e-27, 2.695996e-26, 
    5.269447e-26, 1.225453e-26, -8.578169e-27, -8.087988e-26, 2.818541e-26, 
    9.803622e-26, 1.053889e-25, 9.558531e-26, 7.475262e-26, 3.921449e-26, 
    1.715634e-26, 2.818541e-26, 1.102908e-26, 7.842898e-26, 1.225453e-26, 
    -2.818541e-26, 8.578169e-27, -2.205815e-26, 3.308722e-26, -2.573451e-26, 
    -1.090653e-25, -3.063632e-26, 2.941087e-26,
  1.338114e-32, 1.338112e-32, 1.338113e-32, 1.338112e-32, 1.338112e-32, 
    1.338111e-32, 1.338113e-32, 1.338112e-32, 1.338113e-32, 1.338113e-32, 
    1.338109e-32, 1.338111e-32, 1.338107e-32, 1.338109e-32, 1.338105e-32, 
    1.338107e-32, 1.338105e-32, 1.338105e-32, 1.338104e-32, 1.338104e-32, 
    1.338102e-32, 1.338104e-32, 1.338101e-32, 1.338103e-32, 1.338102e-32, 
    1.338104e-32, 1.338111e-32, 1.33811e-32, 1.338111e-32, 1.338111e-32, 
    1.338111e-32, 1.338112e-32, 1.338113e-32, 1.338114e-32, 1.338113e-32, 
    1.338113e-32, 1.338111e-32, 1.338111e-32, 1.33811e-32, 1.33811e-32, 
    1.338108e-32, 1.338109e-32, 1.338106e-32, 1.338107e-32, 1.338104e-32, 
    1.338105e-32, 1.338104e-32, 1.338104e-32, 1.338104e-32, 1.338105e-32, 
    1.338105e-32, 1.338106e-32, 1.338109e-32, 1.338108e-32, 1.33811e-32, 
    1.338112e-32, 1.338113e-32, 1.338114e-32, 1.338114e-32, 1.338114e-32, 
    1.338113e-32, 1.338112e-32, 1.338111e-32, 1.33811e-32, 1.33811e-32, 
    1.338108e-32, 1.338108e-32, 1.338106e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338104e-32, 1.338104e-32, 1.338105e-32, 
    1.338104e-32, 1.338106e-32, 1.338106e-32, 1.33811e-32, 1.338111e-32, 
    1.338112e-32, 1.338113e-32, 1.338114e-32, 1.338113e-32, 1.338113e-32, 
    1.338112e-32, 1.338112e-32, 1.338112e-32, 1.33811e-32, 1.338111e-32, 
    1.338107e-32, 1.338109e-32, 1.338105e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338105e-32, 1.338104e-32, 1.338103e-32, 
    1.338104e-32, 1.338103e-32, 1.338105e-32, 1.338104e-32, 1.338112e-32, 
    1.338112e-32, 1.338112e-32, 1.338113e-32, 1.338113e-32, 1.338114e-32, 
    1.338113e-32, 1.338113e-32, 1.338112e-32, 1.338111e-32, 1.338111e-32, 
    1.33811e-32, 1.338109e-32, 1.338107e-32, 1.338106e-32, 1.338105e-32, 
    1.338106e-32, 1.338105e-32, 1.338106e-32, 1.338106e-32, 1.338103e-32, 
    1.338105e-32, 1.338103e-32, 1.338103e-32, 1.338104e-32, 1.338103e-32, 
    1.338112e-32, 1.338112e-32, 1.338113e-32, 1.338113e-32, 1.338114e-32, 
    1.338113e-32, 1.338113e-32, 1.338111e-32, 1.338111e-32, 1.33811e-32, 
    1.33811e-32, 1.338109e-32, 1.338107e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 
    1.338104e-32, 1.338105e-32, 1.338103e-32, 1.338103e-32, 1.338103e-32, 
    1.338103e-32, 1.338112e-32, 1.338112e-32, 1.338112e-32, 1.338112e-32, 
    1.338112e-32, 1.33811e-32, 1.33811e-32, 1.338108e-32, 1.338109e-32, 
    1.338108e-32, 1.338109e-32, 1.338109e-32, 1.338108e-32, 1.338109e-32, 
    1.338106e-32, 1.338108e-32, 1.338105e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338104e-32, 1.338103e-32, 1.338102e-32, 
    1.338102e-32, 1.338102e-32, 1.338111e-32, 1.33811e-32, 1.338111e-32, 
    1.33811e-32, 1.338109e-32, 1.338109e-32, 1.338107e-32, 1.338108e-32, 
    1.338107e-32, 1.338106e-32, 1.338108e-32, 1.338107e-32, 1.33811e-32, 
    1.33811e-32, 1.33811e-32, 1.338111e-32, 1.338107e-32, 1.338109e-32, 
    1.338106e-32, 1.338107e-32, 1.338104e-32, 1.338105e-32, 1.338103e-32, 
    1.338101e-32, 1.3381e-32, 1.338099e-32, 1.33811e-32, 1.338111e-32, 
    1.33811e-32, 1.338109e-32, 1.338108e-32, 1.338107e-32, 1.338107e-32, 
    1.338107e-32, 1.338106e-32, 1.338105e-32, 1.338106e-32, 1.338105e-32, 
    1.338109e-32, 1.338107e-32, 1.338111e-32, 1.33811e-32, 1.338109e-32, 
    1.338109e-32, 1.338108e-32, 1.338107e-32, 1.338106e-32, 1.338107e-32, 
    1.338102e-32, 1.338104e-32, 1.338098e-32, 1.338099e-32, 1.338111e-32, 
    1.33811e-32, 1.338108e-32, 1.338109e-32, 1.338107e-32, 1.338106e-32, 
    1.338106e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 
    1.338105e-32, 1.338107e-32, 1.338106e-32, 1.338109e-32, 1.338108e-32, 
    1.338108e-32, 1.338109e-32, 1.338108e-32, 1.338106e-32, 1.338106e-32, 
    1.338106e-32, 1.338105e-32, 1.338107e-32, 1.338101e-32, 1.338105e-32, 
    1.33811e-32, 1.338109e-32, 1.338108e-32, 1.338109e-32, 1.338106e-32, 
    1.338107e-32, 1.338105e-32, 1.338105e-32, 1.338104e-32, 1.338105e-32, 
    1.338105e-32, 1.338105e-32, 1.338106e-32, 1.338107e-32, 1.338108e-32, 
    1.338109e-32, 1.338109e-32, 1.338108e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338107e-32, 1.338106e-32, 1.338106e-32, 
    1.338105e-32, 1.338108e-32, 1.338105e-32, 1.338108e-32, 1.338108e-32, 
    1.338107e-32, 1.338106e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 
    1.338106e-32, 1.338107e-32, 1.338107e-32, 1.338107e-32, 1.338108e-32, 
    1.338108e-32, 1.338108e-32, 1.338108e-32, 1.338106e-32, 1.338105e-32, 
    1.338104e-32, 1.338104e-32, 1.338102e-32, 1.338103e-32, 1.338101e-32, 
    1.338103e-32, 1.3381e-32, 1.338105e-32, 1.338103e-32, 1.338107e-32, 
    1.338107e-32, 1.338106e-32, 1.338104e-32, 1.338105e-32, 1.338104e-32, 
    1.338107e-32, 1.338108e-32, 1.338108e-32, 1.338109e-32, 1.338108e-32, 
    1.338108e-32, 1.338108e-32, 1.338108e-32, 1.338106e-32, 1.338107e-32, 
    1.338105e-32, 1.338104e-32, 1.338102e-32, 1.3381e-32, 1.338099e-32, 
    1.338098e-32, 1.338098e-32, 1.338098e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.70699e-15, 1.711335e-15, 1.710491e-15, 1.713992e-15, 1.712051e-15, 
    1.714342e-15, 1.707872e-15, 1.711507e-15, 1.709187e-15, 1.707382e-15, 
    1.720775e-15, 1.714148e-15, 1.727653e-15, 1.723435e-15, 1.734024e-15, 
    1.726996e-15, 1.73544e-15, 1.733823e-15, 1.738691e-15, 1.737297e-15, 
    1.743512e-15, 1.739334e-15, 1.746732e-15, 1.742516e-15, 1.743175e-15, 
    1.739195e-15, 1.715484e-15, 1.71995e-15, 1.715219e-15, 1.715856e-15, 
    1.715571e-15, 1.71209e-15, 1.710334e-15, 1.706658e-15, 1.707326e-15, 
    1.710026e-15, 1.716143e-15, 1.714069e-15, 1.719297e-15, 1.719179e-15, 
    1.72499e-15, 1.722371e-15, 1.732126e-15, 1.729357e-15, 1.737355e-15, 
    1.735345e-15, 1.73726e-15, 1.73668e-15, 1.737268e-15, 1.73432e-15, 
    1.735583e-15, 1.732988e-15, 1.722862e-15, 1.72584e-15, 1.716949e-15, 
    1.71159e-15, 1.708031e-15, 1.705502e-15, 1.705859e-15, 1.706541e-15, 
    1.710042e-15, 1.713333e-15, 1.715838e-15, 1.717513e-15, 1.719162e-15, 
    1.724147e-15, 1.726786e-15, 1.732685e-15, 1.731623e-15, 1.733423e-15, 
    1.735145e-15, 1.738032e-15, 1.737557e-15, 1.738828e-15, 1.733377e-15, 
    1.737e-15, 1.731017e-15, 1.732654e-15, 1.719605e-15, 1.714629e-15, 
    1.712507e-15, 1.710653e-15, 1.706134e-15, 1.709255e-15, 1.708025e-15, 
    1.710952e-15, 1.71281e-15, 1.711891e-15, 1.717558e-15, 1.715356e-15, 
    1.726942e-15, 1.721956e-15, 1.734944e-15, 1.731841e-15, 1.735688e-15, 
    1.733726e-15, 1.737087e-15, 1.734062e-15, 1.739301e-15, 1.740441e-15, 
    1.739662e-15, 1.742654e-15, 1.733894e-15, 1.73726e-15, 1.711865e-15, 
    1.712015e-15, 1.712713e-15, 1.709642e-15, 1.709455e-15, 1.70664e-15, 
    1.709145e-15, 1.710211e-15, 1.712918e-15, 1.714517e-15, 1.716037e-15, 
    1.719376e-15, 1.723102e-15, 1.728307e-15, 1.732042e-15, 1.734543e-15, 
    1.73301e-15, 1.734364e-15, 1.73285e-15, 1.732141e-15, 1.740013e-15, 
    1.735595e-15, 1.742223e-15, 1.741857e-15, 1.738858e-15, 1.741898e-15, 
    1.71212e-15, 1.711258e-15, 1.708261e-15, 1.710607e-15, 1.706333e-15, 
    1.708725e-15, 1.710099e-15, 1.715401e-15, 1.716566e-15, 1.717644e-15, 
    1.719774e-15, 1.722505e-15, 1.727291e-15, 1.731451e-15, 1.735245e-15, 
    1.734968e-15, 1.735065e-15, 1.735912e-15, 1.733814e-15, 1.736256e-15, 
    1.736666e-15, 1.735595e-15, 1.741808e-15, 1.740034e-15, 1.741849e-15, 
    1.740695e-15, 1.711538e-15, 1.712989e-15, 1.712205e-15, 1.713679e-15, 
    1.71264e-15, 1.717255e-15, 1.718638e-15, 1.725101e-15, 1.722451e-15, 
    1.72667e-15, 1.72288e-15, 1.723552e-15, 1.726805e-15, 1.723086e-15, 
    1.731221e-15, 1.725706e-15, 1.735945e-15, 1.730442e-15, 1.736289e-15, 
    1.735229e-15, 1.736985e-15, 1.738556e-15, 1.740533e-15, 1.744175e-15, 
    1.743332e-15, 1.746377e-15, 1.715152e-15, 1.717031e-15, 1.716866e-15, 
    1.718833e-15, 1.720287e-15, 1.723436e-15, 1.728481e-15, 1.726585e-15, 
    1.730066e-15, 1.730765e-15, 1.725476e-15, 1.728723e-15, 1.718289e-15, 
    1.719976e-15, 1.718972e-15, 1.715299e-15, 1.727021e-15, 1.721009e-15, 
    1.732103e-15, 1.728853e-15, 1.738332e-15, 1.73362e-15, 1.742868e-15, 
    1.746811e-15, 1.750523e-15, 1.754851e-15, 1.718057e-15, 1.716781e-15, 
    1.719067e-15, 1.722226e-15, 1.725158e-15, 1.729051e-15, 1.72945e-15, 
    1.730178e-15, 1.732065e-15, 1.733651e-15, 1.730407e-15, 1.734048e-15, 
    1.720365e-15, 1.727543e-15, 1.716297e-15, 1.719685e-15, 1.722041e-15, 
    1.721009e-15, 1.726369e-15, 1.727631e-15, 1.732753e-15, 1.730107e-15, 
    1.745838e-15, 1.738886e-15, 1.758145e-15, 1.752774e-15, 1.716334e-15, 
    1.718053e-15, 1.724029e-15, 1.721187e-15, 1.729311e-15, 1.731308e-15, 
    1.732931e-15, 1.735003e-15, 1.735227e-15, 1.736454e-15, 1.734443e-15, 
    1.736375e-15, 1.729059e-15, 1.732331e-15, 1.723348e-15, 1.725535e-15, 
    1.72453e-15, 1.723425e-15, 1.726833e-15, 1.730458e-15, 1.730537e-15, 
    1.731699e-15, 1.734966e-15, 1.729344e-15, 1.746731e-15, 1.736001e-15, 
    1.719927e-15, 1.723232e-15, 1.723706e-15, 1.722426e-15, 1.731107e-15, 
    1.727964e-15, 1.736425e-15, 1.73414e-15, 1.737883e-15, 1.736023e-15, 
    1.73575e-15, 1.73336e-15, 1.731872e-15, 1.728108e-15, 1.725043e-15, 
    1.722612e-15, 1.723177e-15, 1.725848e-15, 1.73068e-15, 1.735247e-15, 
    1.734247e-15, 1.737599e-15, 1.728723e-15, 1.732446e-15, 1.731007e-15, 
    1.734759e-15, 1.726535e-15, 1.733534e-15, 1.724743e-15, 1.725515e-15, 
    1.727902e-15, 1.732698e-15, 1.73376e-15, 1.734892e-15, 1.734194e-15, 
    1.730803e-15, 1.730248e-15, 1.727844e-15, 1.727179e-15, 1.725347e-15, 
    1.723828e-15, 1.725215e-15, 1.726671e-15, 1.730805e-15, 1.734526e-15, 
    1.738578e-15, 1.73957e-15, 1.744293e-15, 1.740446e-15, 1.74679e-15, 
    1.741394e-15, 1.750731e-15, 1.733942e-15, 1.741239e-15, 1.728011e-15, 
    1.729439e-15, 1.732018e-15, 1.73793e-15, 1.734741e-15, 1.738471e-15, 
    1.730226e-15, 1.725939e-15, 1.724831e-15, 1.722759e-15, 1.724878e-15, 
    1.724706e-15, 1.726732e-15, 1.726082e-15, 1.730942e-15, 1.728332e-15, 
    1.735742e-15, 1.738442e-15, 1.746058e-15, 1.750717e-15, 1.755456e-15, 
    1.757545e-15, 1.758181e-15, 1.758446e-15 ;

 LITR3N_vr =
  7.663647e-06, 7.66364e-06, 7.663641e-06, 7.663634e-06, 7.663638e-06, 
    7.663634e-06, 7.663645e-06, 7.663639e-06, 7.663643e-06, 7.663646e-06, 
    7.663622e-06, 7.663634e-06, 7.663611e-06, 7.663618e-06, 7.6636e-06, 
    7.663612e-06, 7.663597e-06, 7.6636e-06, 7.663592e-06, 7.663594e-06, 
    7.663583e-06, 7.663591e-06, 7.663578e-06, 7.663585e-06, 7.663583e-06, 
    7.663591e-06, 7.663632e-06, 7.663624e-06, 7.663632e-06, 7.663632e-06, 
    7.663632e-06, 7.663638e-06, 7.663641e-06, 7.663648e-06, 7.663646e-06, 
    7.663642e-06, 7.663631e-06, 7.663634e-06, 7.663625e-06, 7.663626e-06, 
    7.663615e-06, 7.66362e-06, 7.663603e-06, 7.663608e-06, 7.663594e-06, 
    7.663597e-06, 7.663594e-06, 7.663595e-06, 7.663594e-06, 7.663599e-06, 
    7.663597e-06, 7.663602e-06, 7.663619e-06, 7.663614e-06, 7.66363e-06, 
    7.663639e-06, 7.663645e-06, 7.66365e-06, 7.663649e-06, 7.663648e-06, 
    7.663642e-06, 7.663636e-06, 7.663632e-06, 7.663629e-06, 7.663626e-06, 
    7.663617e-06, 7.663612e-06, 7.663602e-06, 7.663604e-06, 7.663601e-06, 
    7.663598e-06, 7.663592e-06, 7.663593e-06, 7.663592e-06, 7.663601e-06, 
    7.663594e-06, 7.663605e-06, 7.663602e-06, 7.663625e-06, 7.663633e-06, 
    7.663637e-06, 7.663641e-06, 7.663649e-06, 7.663643e-06, 7.663645e-06, 
    7.66364e-06, 7.663637e-06, 7.663639e-06, 7.663629e-06, 7.663632e-06, 
    7.663612e-06, 7.663621e-06, 7.663598e-06, 7.663603e-06, 7.663597e-06, 
    7.663601e-06, 7.663594e-06, 7.6636e-06, 7.663591e-06, 7.663589e-06, 
    7.66359e-06, 7.663584e-06, 7.6636e-06, 7.663594e-06, 7.663639e-06, 
    7.663638e-06, 7.663637e-06, 7.663642e-06, 7.663642e-06, 7.663648e-06, 
    7.663643e-06, 7.663642e-06, 7.663637e-06, 7.663633e-06, 7.663632e-06, 
    7.663625e-06, 7.663619e-06, 7.66361e-06, 7.663603e-06, 7.663599e-06, 
    7.663602e-06, 7.663599e-06, 7.663602e-06, 7.663603e-06, 7.663589e-06, 
    7.663597e-06, 7.663585e-06, 7.663586e-06, 7.663592e-06, 7.663586e-06, 
    7.663638e-06, 7.66364e-06, 7.663644e-06, 7.663641e-06, 7.663648e-06, 
    7.663644e-06, 7.663642e-06, 7.663632e-06, 7.663631e-06, 7.663628e-06, 
    7.663624e-06, 7.66362e-06, 7.663612e-06, 7.663604e-06, 7.663598e-06, 
    7.663598e-06, 7.663598e-06, 7.663596e-06, 7.6636e-06, 7.663596e-06, 
    7.663595e-06, 7.663597e-06, 7.663586e-06, 7.663589e-06, 7.663586e-06, 
    7.663588e-06, 7.663639e-06, 7.663636e-06, 7.663638e-06, 7.663635e-06, 
    7.663637e-06, 7.663629e-06, 7.663627e-06, 7.663615e-06, 7.66362e-06, 
    7.663612e-06, 7.663619e-06, 7.663618e-06, 7.663612e-06, 7.663619e-06, 
    7.663604e-06, 7.663614e-06, 7.663596e-06, 7.663606e-06, 7.663596e-06, 
    7.663598e-06, 7.663594e-06, 7.663592e-06, 7.663588e-06, 7.663582e-06, 
    7.663583e-06, 7.663578e-06, 7.663632e-06, 7.66363e-06, 7.66363e-06, 
    7.663626e-06, 7.663623e-06, 7.663618e-06, 7.66361e-06, 7.663612e-06, 
    7.663607e-06, 7.663605e-06, 7.663614e-06, 7.663609e-06, 7.663627e-06, 
    7.663624e-06, 7.663626e-06, 7.663632e-06, 7.663612e-06, 7.663622e-06, 
    7.663603e-06, 7.663609e-06, 7.663592e-06, 7.663601e-06, 7.663584e-06, 
    7.663577e-06, 7.663571e-06, 7.663563e-06, 7.663628e-06, 7.66363e-06, 
    7.663626e-06, 7.663621e-06, 7.663615e-06, 7.663609e-06, 7.663608e-06, 
    7.663606e-06, 7.663603e-06, 7.663601e-06, 7.663606e-06, 7.6636e-06, 
    7.663623e-06, 7.663611e-06, 7.663631e-06, 7.663625e-06, 7.663621e-06, 
    7.663622e-06, 7.663613e-06, 7.663611e-06, 7.663602e-06, 7.663607e-06, 
    7.663579e-06, 7.663592e-06, 7.663558e-06, 7.663567e-06, 7.663631e-06, 
    7.663628e-06, 7.663617e-06, 7.663622e-06, 7.663608e-06, 7.663604e-06, 
    7.663602e-06, 7.663598e-06, 7.663598e-06, 7.663595e-06, 7.663599e-06, 
    7.663595e-06, 7.663609e-06, 7.663602e-06, 7.663618e-06, 7.663614e-06, 
    7.663616e-06, 7.663618e-06, 7.663612e-06, 7.663606e-06, 7.663606e-06, 
    7.663603e-06, 7.663598e-06, 7.663608e-06, 7.663578e-06, 7.663596e-06, 
    7.663624e-06, 7.663619e-06, 7.663618e-06, 7.66362e-06, 7.663605e-06, 
    7.663611e-06, 7.663595e-06, 7.6636e-06, 7.663593e-06, 7.663596e-06, 
    7.663597e-06, 7.663601e-06, 7.663603e-06, 7.66361e-06, 7.663615e-06, 
    7.66362e-06, 7.663619e-06, 7.663614e-06, 7.663605e-06, 7.663598e-06, 
    7.6636e-06, 7.663593e-06, 7.663609e-06, 7.663602e-06, 7.663605e-06, 
    7.663599e-06, 7.663612e-06, 7.663601e-06, 7.663616e-06, 7.663614e-06, 
    7.663611e-06, 7.663602e-06, 7.6636e-06, 7.663598e-06, 7.6636e-06, 
    7.663605e-06, 7.663606e-06, 7.663611e-06, 7.663612e-06, 7.663615e-06, 
    7.663618e-06, 7.663615e-06, 7.663612e-06, 7.663605e-06, 7.663599e-06, 
    7.663592e-06, 7.66359e-06, 7.663582e-06, 7.663589e-06, 7.663577e-06, 
    7.663587e-06, 7.663571e-06, 7.6636e-06, 7.663587e-06, 7.663611e-06, 
    7.663608e-06, 7.663603e-06, 7.663592e-06, 7.663599e-06, 7.663592e-06, 
    7.663606e-06, 7.663614e-06, 7.663616e-06, 7.66362e-06, 7.663616e-06, 
    7.663616e-06, 7.663612e-06, 7.663613e-06, 7.663605e-06, 7.66361e-06, 
    7.663597e-06, 7.663592e-06, 7.663579e-06, 7.663571e-06, 7.663562e-06, 
    7.663559e-06, 7.663558e-06, 7.663557e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  6.167196e-14, 6.182895e-14, 6.179845e-14, 6.192495e-14, 6.185481e-14, 
    6.19376e-14, 6.170383e-14, 6.183515e-14, 6.175134e-14, 6.168614e-14, 
    6.217002e-14, 6.19306e-14, 6.241851e-14, 6.22661e-14, 6.264869e-14, 
    6.239477e-14, 6.269984e-14, 6.264143e-14, 6.281729e-14, 6.276694e-14, 
    6.299149e-14, 6.284052e-14, 6.310782e-14, 6.295549e-14, 6.297931e-14, 
    6.283553e-14, 6.197886e-14, 6.214021e-14, 6.196928e-14, 6.199231e-14, 
    6.198199e-14, 6.185624e-14, 6.17928e-14, 6.165999e-14, 6.168412e-14, 
    6.178168e-14, 6.200266e-14, 6.192772e-14, 6.211662e-14, 6.211236e-14, 
    6.232231e-14, 6.222769e-14, 6.258012e-14, 6.248006e-14, 6.276904e-14, 
    6.269642e-14, 6.276562e-14, 6.274465e-14, 6.276589e-14, 6.265937e-14, 
    6.270502e-14, 6.261127e-14, 6.22454e-14, 6.235302e-14, 6.203178e-14, 
    6.183818e-14, 6.170958e-14, 6.16182e-14, 6.163113e-14, 6.165575e-14, 
    6.178224e-14, 6.190113e-14, 6.199164e-14, 6.205215e-14, 6.211175e-14, 
    6.229183e-14, 6.238717e-14, 6.260032e-14, 6.256193e-14, 6.262699e-14, 
    6.268919e-14, 6.279349e-14, 6.277634e-14, 6.282225e-14, 6.262531e-14, 
    6.275622e-14, 6.254004e-14, 6.25992e-14, 6.212775e-14, 6.194796e-14, 
    6.18713e-14, 6.180431e-14, 6.164106e-14, 6.175381e-14, 6.170937e-14, 
    6.181511e-14, 6.188223e-14, 6.184904e-14, 6.20538e-14, 6.197423e-14, 
    6.239283e-14, 6.221268e-14, 6.268194e-14, 6.256981e-14, 6.270881e-14, 
    6.263791e-14, 6.275935e-14, 6.265006e-14, 6.283936e-14, 6.288051e-14, 
    6.285238e-14, 6.296047e-14, 6.2644e-14, 6.27656e-14, 6.18481e-14, 
    6.185352e-14, 6.187875e-14, 6.17678e-14, 6.176102e-14, 6.165932e-14, 
    6.174983e-14, 6.178834e-14, 6.188614e-14, 6.194391e-14, 6.199883e-14, 
    6.211949e-14, 6.225408e-14, 6.244212e-14, 6.257708e-14, 6.266745e-14, 
    6.261206e-14, 6.266097e-14, 6.260629e-14, 6.258066e-14, 6.286508e-14, 
    6.270543e-14, 6.294493e-14, 6.29317e-14, 6.282334e-14, 6.293319e-14, 
    6.185732e-14, 6.182617e-14, 6.17179e-14, 6.180264e-14, 6.164824e-14, 
    6.173467e-14, 6.178432e-14, 6.197585e-14, 6.201794e-14, 6.20569e-14, 
    6.213386e-14, 6.223253e-14, 6.240544e-14, 6.255574e-14, 6.269282e-14, 
    6.268278e-14, 6.268631e-14, 6.27169e-14, 6.26411e-14, 6.272934e-14, 
    6.274413e-14, 6.270544e-14, 6.292992e-14, 6.286583e-14, 6.293141e-14, 
    6.288969e-14, 6.18363e-14, 6.188872e-14, 6.18604e-14, 6.191364e-14, 
    6.187612e-14, 6.204285e-14, 6.209279e-14, 6.232632e-14, 6.223058e-14, 
    6.238298e-14, 6.224608e-14, 6.227034e-14, 6.238787e-14, 6.22535e-14, 
    6.254742e-14, 6.234815e-14, 6.271809e-14, 6.251928e-14, 6.273053e-14, 
    6.269223e-14, 6.275566e-14, 6.281243e-14, 6.288384e-14, 6.301545e-14, 
    6.298499e-14, 6.3095e-14, 6.196684e-14, 6.203474e-14, 6.20288e-14, 
    6.209985e-14, 6.215236e-14, 6.226616e-14, 6.244844e-14, 6.237994e-14, 
    6.250571e-14, 6.253093e-14, 6.233986e-14, 6.245717e-14, 6.20802e-14, 
    6.214114e-14, 6.210488e-14, 6.197218e-14, 6.239567e-14, 6.217848e-14, 
    6.25793e-14, 6.246186e-14, 6.280433e-14, 6.263409e-14, 6.296821e-14, 
    6.311069e-14, 6.32448e-14, 6.340114e-14, 6.207183e-14, 6.20257e-14, 
    6.210831e-14, 6.222246e-14, 6.232838e-14, 6.246902e-14, 6.248342e-14, 
    6.250973e-14, 6.257792e-14, 6.263521e-14, 6.251802e-14, 6.264957e-14, 
    6.215519e-14, 6.241453e-14, 6.200823e-14, 6.213065e-14, 6.221575e-14, 
    6.217846e-14, 6.237211e-14, 6.24177e-14, 6.260278e-14, 6.250716e-14, 
    6.307551e-14, 6.282436e-14, 6.352017e-14, 6.332609e-14, 6.200957e-14, 
    6.207169e-14, 6.228758e-14, 6.21849e-14, 6.247842e-14, 6.255055e-14, 
    6.260919e-14, 6.268405e-14, 6.269215e-14, 6.273649e-14, 6.266383e-14, 
    6.273364e-14, 6.246932e-14, 6.258751e-14, 6.226296e-14, 6.234201e-14, 
    6.230566e-14, 6.226576e-14, 6.238888e-14, 6.251985e-14, 6.252271e-14, 
    6.256467e-14, 6.268274e-14, 6.247961e-14, 6.310778e-14, 6.27201e-14, 
    6.213937e-14, 6.225879e-14, 6.227592e-14, 6.222966e-14, 6.254332e-14, 
    6.242975e-14, 6.273542e-14, 6.265289e-14, 6.27881e-14, 6.272093e-14, 
    6.271104e-14, 6.262472e-14, 6.257093e-14, 6.243495e-14, 6.232422e-14, 
    6.223638e-14, 6.225681e-14, 6.235329e-14, 6.252788e-14, 6.269287e-14, 
    6.265673e-14, 6.277783e-14, 6.245716e-14, 6.259169e-14, 6.253969e-14, 
    6.267524e-14, 6.23781e-14, 6.2631e-14, 6.231336e-14, 6.234125e-14, 
    6.242749e-14, 6.260077e-14, 6.263916e-14, 6.268003e-14, 6.265482e-14, 
    6.253232e-14, 6.251226e-14, 6.242541e-14, 6.240139e-14, 6.233519e-14, 
    6.228032e-14, 6.233044e-14, 6.238303e-14, 6.253239e-14, 6.266681e-14, 
    6.281323e-14, 6.284905e-14, 6.301972e-14, 6.288072e-14, 6.310992e-14, 
    6.291497e-14, 6.325231e-14, 6.264573e-14, 6.290935e-14, 6.243144e-14, 
    6.248302e-14, 6.257621e-14, 6.278982e-14, 6.26746e-14, 6.280937e-14, 
    6.251148e-14, 6.235659e-14, 6.231655e-14, 6.224171e-14, 6.231826e-14, 
    6.231204e-14, 6.238525e-14, 6.236174e-14, 6.253735e-14, 6.244305e-14, 
    6.271078e-14, 6.280832e-14, 6.308346e-14, 6.325179e-14, 6.3423e-14, 
    6.349848e-14, 6.352145e-14, 6.353105e-14 ;

 LITTERC =
  5.976081e-05, 5.976067e-05, 5.97607e-05, 5.976058e-05, 5.976064e-05, 
    5.976057e-05, 5.976078e-05, 5.976066e-05, 5.976074e-05, 5.97608e-05, 
    5.976036e-05, 5.976058e-05, 5.976013e-05, 5.976027e-05, 5.975992e-05, 
    5.976015e-05, 5.975987e-05, 5.975993e-05, 5.975977e-05, 5.975981e-05, 
    5.975961e-05, 5.975975e-05, 5.97595e-05, 5.975964e-05, 5.975962e-05, 
    5.975975e-05, 5.976053e-05, 5.976039e-05, 5.976054e-05, 5.976052e-05, 
    5.976053e-05, 5.976064e-05, 5.97607e-05, 5.976082e-05, 5.97608e-05, 
    5.976071e-05, 5.976051e-05, 5.976058e-05, 5.97604e-05, 5.976041e-05, 
    5.976022e-05, 5.976031e-05, 5.975998e-05, 5.976007e-05, 5.975981e-05, 
    5.975988e-05, 5.975981e-05, 5.975983e-05, 5.975981e-05, 5.975991e-05, 
    5.975987e-05, 5.975995e-05, 5.976029e-05, 5.976019e-05, 5.976048e-05, 
    5.976066e-05, 5.976078e-05, 5.976086e-05, 5.976085e-05, 5.976083e-05, 
    5.976071e-05, 5.97606e-05, 5.976052e-05, 5.976047e-05, 5.976041e-05, 
    5.976024e-05, 5.976016e-05, 5.975996e-05, 5.976e-05, 5.975994e-05, 
    5.975988e-05, 5.975979e-05, 5.97598e-05, 5.975976e-05, 5.975994e-05, 
    5.975982e-05, 5.976002e-05, 5.975996e-05, 5.97604e-05, 5.976056e-05, 
    5.976063e-05, 5.976069e-05, 5.976084e-05, 5.976074e-05, 5.976078e-05, 
    5.976068e-05, 5.976062e-05, 5.976065e-05, 5.976046e-05, 5.976054e-05, 
    5.976015e-05, 5.976032e-05, 5.975989e-05, 5.975999e-05, 5.975987e-05, 
    5.975993e-05, 5.975982e-05, 5.975992e-05, 5.975975e-05, 5.975971e-05, 
    5.975974e-05, 5.975964e-05, 5.975992e-05, 5.975981e-05, 5.976065e-05, 
    5.976065e-05, 5.976062e-05, 5.976072e-05, 5.976073e-05, 5.976082e-05, 
    5.976074e-05, 5.976071e-05, 5.976062e-05, 5.976056e-05, 5.976051e-05, 
    5.97604e-05, 5.976028e-05, 5.976011e-05, 5.975999e-05, 5.97599e-05, 
    5.975995e-05, 5.975991e-05, 5.975996e-05, 5.975998e-05, 5.975972e-05, 
    5.975987e-05, 5.975965e-05, 5.975966e-05, 5.975976e-05, 5.975966e-05, 
    5.976064e-05, 5.976067e-05, 5.976077e-05, 5.976069e-05, 5.976083e-05, 
    5.976075e-05, 5.976071e-05, 5.976054e-05, 5.97605e-05, 5.976046e-05, 
    5.976039e-05, 5.97603e-05, 5.976014e-05, 5.976e-05, 5.975988e-05, 
    5.975989e-05, 5.975988e-05, 5.975986e-05, 5.975993e-05, 5.975985e-05, 
    5.975983e-05, 5.975987e-05, 5.975966e-05, 5.975972e-05, 5.975966e-05, 
    5.97597e-05, 5.976066e-05, 5.976062e-05, 5.976064e-05, 5.976059e-05, 
    5.976063e-05, 5.976047e-05, 5.976043e-05, 5.976022e-05, 5.97603e-05, 
    5.976016e-05, 5.976029e-05, 5.976027e-05, 5.976016e-05, 5.976028e-05, 
    5.976001e-05, 5.976019e-05, 5.975986e-05, 5.976004e-05, 5.975984e-05, 
    5.975988e-05, 5.975982e-05, 5.975977e-05, 5.975971e-05, 5.975959e-05, 
    5.975961e-05, 5.975951e-05, 5.976054e-05, 5.976048e-05, 5.976049e-05, 
    5.976042e-05, 5.976037e-05, 5.976027e-05, 5.97601e-05, 5.976016e-05, 
    5.976005e-05, 5.976003e-05, 5.97602e-05, 5.97601e-05, 5.976044e-05, 
    5.976038e-05, 5.976042e-05, 5.976054e-05, 5.976015e-05, 5.976035e-05, 
    5.975998e-05, 5.976009e-05, 5.975978e-05, 5.975994e-05, 5.975963e-05, 
    5.97595e-05, 5.975938e-05, 5.975923e-05, 5.976045e-05, 5.976049e-05, 
    5.976042e-05, 5.976031e-05, 5.976021e-05, 5.976008e-05, 5.976007e-05, 
    5.976005e-05, 5.975999e-05, 5.975993e-05, 5.976004e-05, 5.975992e-05, 
    5.976037e-05, 5.976014e-05, 5.976051e-05, 5.976039e-05, 5.976032e-05, 
    5.976035e-05, 5.976017e-05, 5.976013e-05, 5.975996e-05, 5.976005e-05, 
    5.975953e-05, 5.975976e-05, 5.975912e-05, 5.97593e-05, 5.97605e-05, 
    5.976045e-05, 5.976025e-05, 5.976034e-05, 5.976008e-05, 5.976001e-05, 
    5.975996e-05, 5.975989e-05, 5.975988e-05, 5.975984e-05, 5.975991e-05, 
    5.975984e-05, 5.976008e-05, 5.975998e-05, 5.976027e-05, 5.97602e-05, 
    5.976023e-05, 5.976027e-05, 5.976016e-05, 5.976004e-05, 5.976003e-05, 
    5.976e-05, 5.975989e-05, 5.976007e-05, 5.97595e-05, 5.975986e-05, 
    5.976039e-05, 5.976028e-05, 5.976026e-05, 5.97603e-05, 5.976002e-05, 
    5.976012e-05, 5.975984e-05, 5.975992e-05, 5.975979e-05, 5.975986e-05, 
    5.975986e-05, 5.975994e-05, 5.975999e-05, 5.976012e-05, 5.976022e-05, 
    5.97603e-05, 5.976028e-05, 5.976019e-05, 5.976003e-05, 5.975988e-05, 
    5.975991e-05, 5.97598e-05, 5.97601e-05, 5.975997e-05, 5.976002e-05, 
    5.97599e-05, 5.976017e-05, 5.975994e-05, 5.976023e-05, 5.97602e-05, 
    5.976012e-05, 5.975996e-05, 5.975993e-05, 5.975989e-05, 5.975991e-05, 
    5.976003e-05, 5.976004e-05, 5.976012e-05, 5.976015e-05, 5.976021e-05, 
    5.976026e-05, 5.976021e-05, 5.976016e-05, 5.976003e-05, 5.97599e-05, 
    5.975977e-05, 5.975974e-05, 5.975958e-05, 5.975971e-05, 5.97595e-05, 
    5.975968e-05, 5.975937e-05, 5.975992e-05, 5.975968e-05, 5.976012e-05, 
    5.976007e-05, 5.975999e-05, 5.975979e-05, 5.97599e-05, 5.975978e-05, 
    5.976004e-05, 5.976019e-05, 5.976022e-05, 5.976029e-05, 5.976022e-05, 
    5.976023e-05, 5.976016e-05, 5.976018e-05, 5.976002e-05, 5.976011e-05, 
    5.975986e-05, 5.975978e-05, 5.975952e-05, 5.975937e-05, 5.975921e-05, 
    5.975914e-05, 5.975912e-05, 5.975911e-05 ;

 LITTERC_HR =
  9.949716e-13, 9.975021e-13, 9.970106e-13, 9.990496e-13, 9.979191e-13, 
    9.992536e-13, 9.954853e-13, 9.976022e-13, 9.962513e-13, 9.952001e-13, 
    1.003e-12, 9.991407e-13, 1.007005e-12, 1.004549e-12, 1.010716e-12, 
    1.006623e-12, 1.01154e-12, 1.010599e-12, 1.013433e-12, 1.012622e-12, 
    1.016241e-12, 1.013808e-12, 1.018117e-12, 1.015661e-12, 1.016045e-12, 
    1.013728e-12, 9.999188e-13, 1.00252e-12, 9.997643e-13, 1.000136e-12, 
    9.999692e-13, 9.979422e-13, 9.969193e-13, 9.947787e-13, 9.951677e-13, 
    9.967402e-13, 1.000302e-12, 9.990944e-13, 1.002139e-12, 1.002071e-12, 
    1.005455e-12, 1.00393e-12, 1.009611e-12, 1.007998e-12, 1.012656e-12, 
    1.011485e-12, 1.012601e-12, 1.012263e-12, 1.012605e-12, 1.010888e-12, 
    1.011624e-12, 1.010113e-12, 1.004215e-12, 1.00595e-12, 1.000772e-12, 
    9.97651e-13, 9.955781e-13, 9.941052e-13, 9.943135e-13, 9.947103e-13, 
    9.967493e-13, 9.986657e-13, 1.000125e-12, 1.0011e-12, 1.002061e-12, 
    1.004964e-12, 1.0065e-12, 1.009936e-12, 1.009317e-12, 1.010366e-12, 
    1.011369e-12, 1.01305e-12, 1.012773e-12, 1.013513e-12, 1.010339e-12, 
    1.012449e-12, 1.008965e-12, 1.009918e-12, 1.002319e-12, 9.994205e-13, 
    9.981848e-13, 9.971051e-13, 9.944735e-13, 9.962909e-13, 9.955746e-13, 
    9.972791e-13, 9.983611e-13, 9.978262e-13, 1.001127e-12, 9.99844e-13, 
    1.006592e-12, 1.003688e-12, 1.011252e-12, 1.009444e-12, 1.011685e-12, 
    1.010542e-12, 1.0125e-12, 1.010738e-12, 1.013789e-12, 1.014453e-12, 
    1.013999e-12, 1.015741e-12, 1.01064e-12, 1.0126e-12, 9.97811e-13, 
    9.978983e-13, 9.98305e-13, 9.965165e-13, 9.964073e-13, 9.947679e-13, 
    9.96227e-13, 9.968477e-13, 9.98424e-13, 9.993553e-13, 1.00024e-12, 
    1.002185e-12, 1.004355e-12, 1.007386e-12, 1.009562e-12, 1.011018e-12, 
    1.010125e-12, 1.010914e-12, 1.010032e-12, 1.009619e-12, 1.014204e-12, 
    1.01163e-12, 1.015491e-12, 1.015278e-12, 1.013531e-12, 1.015302e-12, 
    9.979595e-13, 9.974574e-13, 9.957122e-13, 9.970781e-13, 9.945893e-13, 
    9.959824e-13, 9.967827e-13, 9.998701e-13, 1.000549e-12, 1.001177e-12, 
    1.002417e-12, 1.004008e-12, 1.006795e-12, 1.009218e-12, 1.011427e-12, 
    1.011265e-12, 1.011322e-12, 1.011815e-12, 1.010594e-12, 1.012016e-12, 
    1.012254e-12, 1.011631e-12, 1.015249e-12, 1.014216e-12, 1.015273e-12, 
    1.014601e-12, 9.976207e-13, 9.984656e-13, 9.980091e-13, 9.988674e-13, 
    9.982625e-13, 1.00095e-12, 1.001755e-12, 1.00552e-12, 1.003976e-12, 
    1.006433e-12, 1.004226e-12, 1.004617e-12, 1.006512e-12, 1.004346e-12, 
    1.009083e-12, 1.005871e-12, 1.011834e-12, 1.00863e-12, 1.012035e-12, 
    1.011418e-12, 1.01244e-12, 1.013355e-12, 1.014506e-12, 1.016628e-12, 
    1.016137e-12, 1.01791e-12, 9.997249e-13, 1.000819e-12, 1.000724e-12, 
    1.001869e-12, 1.002715e-12, 1.00455e-12, 1.007488e-12, 1.006384e-12, 
    1.008411e-12, 1.008818e-12, 1.005738e-12, 1.007629e-12, 1.001552e-12, 
    1.002534e-12, 1.00195e-12, 9.99811e-13, 1.006637e-12, 1.003136e-12, 
    1.009597e-12, 1.007704e-12, 1.013225e-12, 1.01048e-12, 1.015866e-12, 
    1.018163e-12, 1.020324e-12, 1.022845e-12, 1.001417e-12, 1.000674e-12, 
    1.002005e-12, 1.003845e-12, 1.005553e-12, 1.00782e-12, 1.008052e-12, 
    1.008476e-12, 1.009575e-12, 1.010498e-12, 1.00861e-12, 1.01073e-12, 
    1.002761e-12, 1.006941e-12, 1.000392e-12, 1.002366e-12, 1.003737e-12, 
    1.003136e-12, 1.006258e-12, 1.006993e-12, 1.009976e-12, 1.008434e-12, 
    1.017596e-12, 1.013548e-12, 1.024763e-12, 1.021635e-12, 1.000414e-12, 
    1.001415e-12, 1.004895e-12, 1.00324e-12, 1.007971e-12, 1.009134e-12, 
    1.010079e-12, 1.011286e-12, 1.011416e-12, 1.012131e-12, 1.01096e-12, 
    1.012085e-12, 1.007824e-12, 1.00973e-12, 1.004498e-12, 1.005772e-12, 
    1.005186e-12, 1.004543e-12, 1.006528e-12, 1.008639e-12, 1.008685e-12, 
    1.009362e-12, 1.011265e-12, 1.00799e-12, 1.018116e-12, 1.011867e-12, 
    1.002506e-12, 1.004431e-12, 1.004707e-12, 1.003961e-12, 1.009017e-12, 
    1.007187e-12, 1.012114e-12, 1.010784e-12, 1.012963e-12, 1.01188e-12, 
    1.011721e-12, 1.010329e-12, 1.009462e-12, 1.00727e-12, 1.005486e-12, 
    1.00407e-12, 1.004399e-12, 1.005954e-12, 1.008768e-12, 1.011428e-12, 
    1.010845e-12, 1.012797e-12, 1.007628e-12, 1.009797e-12, 1.008959e-12, 
    1.011144e-12, 1.006354e-12, 1.010431e-12, 1.005311e-12, 1.00576e-12, 
    1.00715e-12, 1.009943e-12, 1.010562e-12, 1.011221e-12, 1.010815e-12, 
    1.00884e-12, 1.008517e-12, 1.007117e-12, 1.00673e-12, 1.005662e-12, 
    1.004778e-12, 1.005586e-12, 1.006434e-12, 1.008841e-12, 1.011008e-12, 
    1.013368e-12, 1.013946e-12, 1.016696e-12, 1.014456e-12, 1.01815e-12, 
    1.015008e-12, 1.020446e-12, 1.010668e-12, 1.014917e-12, 1.007214e-12, 
    1.008045e-12, 1.009548e-12, 1.012991e-12, 1.011134e-12, 1.013306e-12, 
    1.008504e-12, 1.006007e-12, 1.005362e-12, 1.004156e-12, 1.00539e-12, 
    1.005289e-12, 1.006469e-12, 1.00609e-12, 1.008921e-12, 1.007401e-12, 
    1.011717e-12, 1.013289e-12, 1.017724e-12, 1.020437e-12, 1.023197e-12, 
    1.024414e-12, 1.024784e-12, 1.024938e-12 ;

 LITTERC_LOSS =
  1.842679e-12, 1.847365e-12, 1.846455e-12, 1.850231e-12, 1.848137e-12, 
    1.850609e-12, 1.84363e-12, 1.847551e-12, 1.845049e-12, 1.843102e-12, 
    1.857547e-12, 1.8504e-12, 1.864965e-12, 1.860416e-12, 1.871837e-12, 
    1.864257e-12, 1.873364e-12, 1.87162e-12, 1.87687e-12, 1.875367e-12, 
    1.882071e-12, 1.877564e-12, 1.885544e-12, 1.880996e-12, 1.881707e-12, 
    1.877415e-12, 1.851841e-12, 1.856658e-12, 1.851555e-12, 1.852242e-12, 
    1.851934e-12, 1.84818e-12, 1.846286e-12, 1.842321e-12, 1.843042e-12, 
    1.845954e-12, 1.852551e-12, 1.850314e-12, 1.855953e-12, 1.855826e-12, 
    1.862094e-12, 1.859269e-12, 1.86979e-12, 1.866803e-12, 1.87543e-12, 
    1.873262e-12, 1.875328e-12, 1.874702e-12, 1.875336e-12, 1.872156e-12, 
    1.873519e-12, 1.87072e-12, 1.859798e-12, 1.86301e-12, 1.853421e-12, 
    1.847641e-12, 1.843802e-12, 1.841074e-12, 1.841459e-12, 1.842195e-12, 
    1.845971e-12, 1.84952e-12, 1.852222e-12, 1.854028e-12, 1.855808e-12, 
    1.861184e-12, 1.86403e-12, 1.870393e-12, 1.869247e-12, 1.871189e-12, 
    1.873046e-12, 1.87616e-12, 1.875648e-12, 1.877019e-12, 1.871139e-12, 
    1.875047e-12, 1.868594e-12, 1.87036e-12, 1.856286e-12, 1.850918e-12, 
    1.84863e-12, 1.84663e-12, 1.841756e-12, 1.845122e-12, 1.843795e-12, 
    1.846952e-12, 1.848956e-12, 1.847965e-12, 1.854078e-12, 1.851702e-12, 
    1.864199e-12, 1.858821e-12, 1.87283e-12, 1.869482e-12, 1.873632e-12, 
    1.871515e-12, 1.875141e-12, 1.871878e-12, 1.877529e-12, 1.878758e-12, 
    1.877918e-12, 1.881145e-12, 1.871697e-12, 1.875327e-12, 1.847937e-12, 
    1.848099e-12, 1.848852e-12, 1.84554e-12, 1.845337e-12, 1.842301e-12, 
    1.845004e-12, 1.846153e-12, 1.849073e-12, 1.850797e-12, 1.852437e-12, 
    1.856039e-12, 1.860057e-12, 1.86567e-12, 1.869699e-12, 1.872397e-12, 
    1.870744e-12, 1.872204e-12, 1.870571e-12, 1.869806e-12, 1.878297e-12, 
    1.873531e-12, 1.880681e-12, 1.880286e-12, 1.877051e-12, 1.88033e-12, 
    1.848212e-12, 1.847282e-12, 1.84405e-12, 1.84658e-12, 1.841971e-12, 
    1.844551e-12, 1.846033e-12, 1.851751e-12, 1.853007e-12, 1.85417e-12, 
    1.856468e-12, 1.859413e-12, 1.864576e-12, 1.869062e-12, 1.873155e-12, 
    1.872855e-12, 1.87296e-12, 1.873873e-12, 1.871611e-12, 1.874245e-12, 
    1.874686e-12, 1.873531e-12, 1.880233e-12, 1.878319e-12, 1.880277e-12, 
    1.879032e-12, 1.847585e-12, 1.84915e-12, 1.848304e-12, 1.849894e-12, 
    1.848773e-12, 1.853751e-12, 1.855242e-12, 1.862214e-12, 1.859355e-12, 
    1.863905e-12, 1.859818e-12, 1.860542e-12, 1.864051e-12, 1.860039e-12, 
    1.868814e-12, 1.862865e-12, 1.873909e-12, 1.867974e-12, 1.87428e-12, 
    1.873137e-12, 1.875031e-12, 1.876725e-12, 1.878857e-12, 1.882786e-12, 
    1.881877e-12, 1.885161e-12, 1.851482e-12, 1.853509e-12, 1.853332e-12, 
    1.855453e-12, 1.85702e-12, 1.860418e-12, 1.865859e-12, 1.863814e-12, 
    1.867569e-12, 1.868322e-12, 1.862618e-12, 1.86612e-12, 1.854866e-12, 
    1.856685e-12, 1.855603e-12, 1.851641e-12, 1.864284e-12, 1.8578e-12, 
    1.869766e-12, 1.86626e-12, 1.876483e-12, 1.871401e-12, 1.881376e-12, 
    1.885629e-12, 1.889633e-12, 1.8943e-12, 1.854616e-12, 1.853239e-12, 
    1.855705e-12, 1.859113e-12, 1.862275e-12, 1.866473e-12, 1.866903e-12, 
    1.867689e-12, 1.869724e-12, 1.871435e-12, 1.867936e-12, 1.871863e-12, 
    1.857105e-12, 1.864847e-12, 1.852717e-12, 1.856372e-12, 1.858913e-12, 
    1.857799e-12, 1.86358e-12, 1.864942e-12, 1.870467e-12, 1.867612e-12, 
    1.884579e-12, 1.877081e-12, 1.897853e-12, 1.892059e-12, 1.852758e-12, 
    1.854612e-12, 1.861057e-12, 1.857992e-12, 1.866754e-12, 1.868907e-12, 
    1.870658e-12, 1.872893e-12, 1.873135e-12, 1.874458e-12, 1.872289e-12, 
    1.874373e-12, 1.866482e-12, 1.870011e-12, 1.860322e-12, 1.862682e-12, 
    1.861597e-12, 1.860405e-12, 1.864081e-12, 1.867991e-12, 1.868076e-12, 
    1.869329e-12, 1.872853e-12, 1.866789e-12, 1.885542e-12, 1.873969e-12, 
    1.856633e-12, 1.860198e-12, 1.860709e-12, 1.859328e-12, 1.868691e-12, 
    1.865301e-12, 1.874426e-12, 1.871963e-12, 1.875999e-12, 1.873994e-12, 
    1.873698e-12, 1.871122e-12, 1.869516e-12, 1.865456e-12, 1.862151e-12, 
    1.859528e-12, 1.860138e-12, 1.863018e-12, 1.86823e-12, 1.873156e-12, 
    1.872077e-12, 1.875693e-12, 1.866119e-12, 1.870136e-12, 1.868583e-12, 
    1.87263e-12, 1.863759e-12, 1.871309e-12, 1.861826e-12, 1.862659e-12, 
    1.865234e-12, 1.870407e-12, 1.871553e-12, 1.872773e-12, 1.87202e-12, 
    1.868363e-12, 1.867764e-12, 1.865172e-12, 1.864455e-12, 1.862478e-12, 
    1.86084e-12, 1.862336e-12, 1.863907e-12, 1.868365e-12, 1.872378e-12, 
    1.876749e-12, 1.877819e-12, 1.882913e-12, 1.878764e-12, 1.885606e-12, 
    1.879786e-12, 1.889857e-12, 1.871749e-12, 1.879618e-12, 1.865351e-12, 
    1.866891e-12, 1.869673e-12, 1.87605e-12, 1.872611e-12, 1.876634e-12, 
    1.867741e-12, 1.863117e-12, 1.861922e-12, 1.859688e-12, 1.861973e-12, 
    1.861787e-12, 1.863973e-12, 1.863271e-12, 1.868513e-12, 1.865698e-12, 
    1.87369e-12, 1.876603e-12, 1.884816e-12, 1.889841e-12, 1.894953e-12, 
    1.897206e-12, 1.897891e-12, 1.898178e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.71279e-18, 1.713045e-18, 1.712998e-18, 1.713193e-18, 1.713087e-18, 
    1.713213e-18, 1.712842e-18, 1.713052e-18, 1.712916e-18, 1.712816e-18, 
    1.713565e-18, 1.713203e-18, 1.713965e-18, 1.713729e-18, 1.714329e-18, 
    1.713926e-18, 1.714411e-18, 1.714323e-18, 1.714603e-18, 1.714523e-18, 
    1.71487e-18, 1.71464e-18, 1.71506e-18, 1.714818e-18, 1.714854e-18, 
    1.714631e-18, 1.713281e-18, 1.713518e-18, 1.713265e-18, 1.713299e-18, 
    1.713285e-18, 1.713087e-18, 1.712984e-18, 1.712775e-18, 1.712812e-18, 
    1.71297e-18, 1.713315e-18, 1.713201e-18, 1.713498e-18, 1.713491e-18, 
    1.713818e-18, 1.713671e-18, 1.714226e-18, 1.714069e-18, 1.714526e-18, 
    1.71441e-18, 1.71452e-18, 1.714487e-18, 1.71452e-18, 1.714351e-18, 
    1.714423e-18, 1.714276e-18, 1.713697e-18, 1.713866e-18, 1.713362e-18, 
    1.713052e-18, 1.71285e-18, 1.71271e-18, 1.71273e-18, 1.712766e-18, 
    1.712971e-18, 1.71316e-18, 1.713302e-18, 1.713396e-18, 1.71349e-18, 
    1.713761e-18, 1.713916e-18, 1.714255e-18, 1.714198e-18, 1.714297e-18, 
    1.714399e-18, 1.714564e-18, 1.714537e-18, 1.714609e-18, 1.714298e-18, 
    1.714503e-18, 1.714165e-18, 1.714257e-18, 1.713498e-18, 1.713233e-18, 
    1.713105e-18, 1.713007e-18, 1.712744e-18, 1.712918e-18, 1.712849e-18, 
    1.713026e-18, 1.71313e-18, 1.713079e-18, 1.713399e-18, 1.713274e-18, 
    1.713925e-18, 1.713644e-18, 1.714387e-18, 1.71421e-18, 1.71443e-18, 
    1.714319e-18, 1.714509e-18, 1.714338e-18, 1.714637e-18, 1.7147e-18, 
    1.714656e-18, 1.714829e-18, 1.714328e-18, 1.714518e-18, 1.713077e-18, 
    1.713085e-18, 1.713125e-18, 1.712949e-18, 1.71293e-18, 1.712773e-18, 
    1.712914e-18, 1.712982e-18, 1.713138e-18, 1.713226e-18, 1.713312e-18, 
    1.713501e-18, 1.713709e-18, 1.714005e-18, 1.714221e-18, 1.714365e-18, 
    1.714278e-18, 1.714355e-18, 1.714269e-18, 1.714229e-18, 1.714675e-18, 
    1.714423e-18, 1.714804e-18, 1.714784e-18, 1.71461e-18, 1.714786e-18, 
    1.713091e-18, 1.713044e-18, 1.712864e-18, 1.713007e-18, 1.712757e-18, 
    1.712889e-18, 1.712973e-18, 1.713273e-18, 1.713343e-18, 1.713402e-18, 
    1.713524e-18, 1.713678e-18, 1.713948e-18, 1.714186e-18, 1.714406e-18, 
    1.71439e-18, 1.714395e-18, 1.714443e-18, 1.714323e-18, 1.714462e-18, 
    1.714484e-18, 1.714425e-18, 1.714781e-18, 1.714679e-18, 1.714783e-18, 
    1.714718e-18, 1.71306e-18, 1.71314e-18, 1.713097e-18, 1.713178e-18, 
    1.713119e-18, 1.713376e-18, 1.713454e-18, 1.71382e-18, 1.713674e-18, 
    1.713912e-18, 1.7137e-18, 1.713736e-18, 1.713912e-18, 1.713712e-18, 
    1.714169e-18, 1.713853e-18, 1.714444e-18, 1.714121e-18, 1.714464e-18, 
    1.714405e-18, 1.714505e-18, 1.714593e-18, 1.714708e-18, 1.714914e-18, 
    1.714867e-18, 1.715042e-18, 1.713263e-18, 1.713366e-18, 1.71336e-18, 
    1.713471e-18, 1.713552e-18, 1.713732e-18, 1.714017e-18, 1.713911e-18, 
    1.71411e-18, 1.714149e-18, 1.713849e-18, 1.71403e-18, 1.713438e-18, 
    1.71353e-18, 1.713477e-18, 1.713269e-18, 1.713931e-18, 1.713589e-18, 
    1.714224e-18, 1.714039e-18, 1.71458e-18, 1.714308e-18, 1.71484e-18, 
    1.715059e-18, 1.715282e-18, 1.715524e-18, 1.713426e-18, 1.713356e-18, 
    1.713485e-18, 1.713658e-18, 1.713829e-18, 1.71405e-18, 1.714075e-18, 
    1.714115e-18, 1.714224e-18, 1.714314e-18, 1.714125e-18, 1.714337e-18, 
    1.713544e-18, 1.713962e-18, 1.713326e-18, 1.713512e-18, 1.713649e-18, 
    1.713593e-18, 1.7139e-18, 1.713971e-18, 1.714259e-18, 1.714112e-18, 
    1.715002e-18, 1.714607e-18, 1.71572e-18, 1.715406e-18, 1.71333e-18, 
    1.713428e-18, 1.713762e-18, 1.713603e-18, 1.714067e-18, 1.714179e-18, 
    1.714274e-18, 1.714389e-18, 1.714404e-18, 1.714473e-18, 1.71436e-18, 
    1.71447e-18, 1.71405e-18, 1.714238e-18, 1.713728e-18, 1.71385e-18, 
    1.713795e-18, 1.713732e-18, 1.713926e-18, 1.714127e-18, 1.714136e-18, 
    1.7142e-18, 1.714369e-18, 1.714069e-18, 1.715043e-18, 1.714431e-18, 
    1.713533e-18, 1.713714e-18, 1.713746e-18, 1.713675e-18, 1.714168e-18, 
    1.713989e-18, 1.714472e-18, 1.714342e-18, 1.714556e-18, 1.714449e-18, 
    1.714433e-18, 1.714298e-18, 1.714212e-18, 1.713996e-18, 1.713821e-18, 
    1.713686e-18, 1.713718e-18, 1.713867e-18, 1.71414e-18, 1.714403e-18, 
    1.714345e-18, 1.71454e-18, 1.714033e-18, 1.714242e-18, 1.71416e-18, 
    1.714377e-18, 1.713907e-18, 1.71429e-18, 1.713807e-18, 1.713851e-18, 
    1.713985e-18, 1.714253e-18, 1.714321e-18, 1.714383e-18, 1.714345e-18, 
    1.714148e-18, 1.714118e-18, 1.713983e-18, 1.713943e-18, 1.713842e-18, 
    1.713755e-18, 1.713833e-18, 1.713913e-18, 1.71415e-18, 1.714361e-18, 
    1.714594e-18, 1.714653e-18, 1.714911e-18, 1.714693e-18, 1.715045e-18, 
    1.714735e-18, 1.715279e-18, 1.714321e-18, 1.714737e-18, 1.713993e-18, 
    1.714074e-18, 1.714215e-18, 1.714552e-18, 1.714376e-18, 1.714584e-18, 
    1.714118e-18, 1.713869e-18, 1.713812e-18, 1.713693e-18, 1.713814e-18, 
    1.713805e-18, 1.713921e-18, 1.713884e-18, 1.714159e-18, 1.714011e-18, 
    1.714432e-18, 1.714584e-18, 1.715021e-18, 1.715287e-18, 1.715566e-18, 
    1.715687e-18, 1.715724e-18, 1.71574e-18 ;

 MEG_acetic_acid =
  2.569186e-19, 2.569567e-19, 2.569497e-19, 2.56979e-19, 2.56963e-19, 
    2.56982e-19, 2.569264e-19, 2.569578e-19, 2.569374e-19, 2.569223e-19, 
    2.570348e-19, 2.569804e-19, 2.570948e-19, 2.570594e-19, 2.571493e-19, 
    2.570888e-19, 2.571617e-19, 2.571484e-19, 2.571904e-19, 2.571784e-19, 
    2.572305e-19, 2.57196e-19, 2.572589e-19, 2.572227e-19, 2.572281e-19, 
    2.571947e-19, 2.569921e-19, 2.570277e-19, 2.569898e-19, 2.569949e-19, 
    2.569928e-19, 2.569631e-19, 2.569476e-19, 2.569163e-19, 2.569219e-19, 
    2.569456e-19, 2.569972e-19, 2.569802e-19, 2.570247e-19, 2.570237e-19, 
    2.570727e-19, 2.570506e-19, 2.571338e-19, 2.571104e-19, 2.571789e-19, 
    2.571615e-19, 2.57178e-19, 2.571731e-19, 2.57178e-19, 2.571526e-19, 
    2.571634e-19, 2.571413e-19, 2.570546e-19, 2.570799e-19, 2.570043e-19, 
    2.569578e-19, 2.569275e-19, 2.569065e-19, 2.569094e-19, 2.56915e-19, 
    2.569457e-19, 2.56974e-19, 2.569953e-19, 2.570095e-19, 2.570236e-19, 
    2.570641e-19, 2.570874e-19, 2.571382e-19, 2.571297e-19, 2.571446e-19, 
    2.571599e-19, 2.571845e-19, 2.571806e-19, 2.571913e-19, 2.571447e-19, 
    2.571754e-19, 2.571247e-19, 2.571385e-19, 2.570246e-19, 2.569849e-19, 
    2.569657e-19, 2.56951e-19, 2.569117e-19, 2.569377e-19, 2.569274e-19, 
    2.569539e-19, 2.569695e-19, 2.569619e-19, 2.570099e-19, 2.569911e-19, 
    2.570888e-19, 2.570467e-19, 2.571581e-19, 2.571315e-19, 2.571645e-19, 
    2.571478e-19, 2.571763e-19, 2.571507e-19, 2.571955e-19, 2.572049e-19, 
    2.571984e-19, 2.572244e-19, 2.571492e-19, 2.571777e-19, 2.569616e-19, 
    2.569628e-19, 2.569688e-19, 2.569423e-19, 2.569394e-19, 2.56916e-19, 
    2.569371e-19, 2.569473e-19, 2.569706e-19, 2.569839e-19, 2.569968e-19, 
    2.570251e-19, 2.570563e-19, 2.571008e-19, 2.571332e-19, 2.571548e-19, 
    2.571417e-19, 2.571533e-19, 2.571403e-19, 2.571343e-19, 2.572012e-19, 
    2.571634e-19, 2.572207e-19, 2.572176e-19, 2.571914e-19, 2.572179e-19, 
    2.569637e-19, 2.569565e-19, 2.569296e-19, 2.56951e-19, 2.569135e-19, 
    2.569334e-19, 2.56946e-19, 2.569909e-19, 2.570014e-19, 2.570103e-19, 
    2.570286e-19, 2.570517e-19, 2.570922e-19, 2.571279e-19, 2.571608e-19, 
    2.571585e-19, 2.571593e-19, 2.571664e-19, 2.571485e-19, 2.571693e-19, 
    2.571726e-19, 2.571637e-19, 2.572171e-19, 2.572019e-19, 2.572175e-19, 
    2.572076e-19, 2.56959e-19, 2.569711e-19, 2.569645e-19, 2.569767e-19, 
    2.569679e-19, 2.570065e-19, 2.57018e-19, 2.57073e-19, 2.570511e-19, 
    2.570868e-19, 2.570549e-19, 2.570604e-19, 2.570868e-19, 2.570568e-19, 
    2.571254e-19, 2.570779e-19, 2.571667e-19, 2.571181e-19, 2.571697e-19, 
    2.571607e-19, 2.571758e-19, 2.57189e-19, 2.572062e-19, 2.57237e-19, 
    2.5723e-19, 2.572563e-19, 2.569894e-19, 2.570049e-19, 2.57004e-19, 
    2.570206e-19, 2.570328e-19, 2.570598e-19, 2.571026e-19, 2.570867e-19, 
    2.571165e-19, 2.571223e-19, 2.570773e-19, 2.571044e-19, 2.570156e-19, 
    2.570294e-19, 2.570216e-19, 2.569903e-19, 2.570896e-19, 2.570383e-19, 
    2.571336e-19, 2.571059e-19, 2.57187e-19, 2.571461e-19, 2.57226e-19, 
    2.572589e-19, 2.572923e-19, 2.573285e-19, 2.570139e-19, 2.570033e-19, 
    2.570227e-19, 2.570487e-19, 2.570743e-19, 2.571075e-19, 2.571112e-19, 
    2.571172e-19, 2.571336e-19, 2.571471e-19, 2.571187e-19, 2.571506e-19, 
    2.570316e-19, 2.570943e-19, 2.569988e-19, 2.570269e-19, 2.570474e-19, 
    2.570389e-19, 2.57085e-19, 2.570957e-19, 2.571389e-19, 2.571168e-19, 
    2.572503e-19, 2.571911e-19, 2.573579e-19, 2.573108e-19, 2.569995e-19, 
    2.570141e-19, 2.570643e-19, 2.570405e-19, 2.5711e-19, 2.571269e-19, 
    2.571411e-19, 2.571584e-19, 2.571606e-19, 2.571709e-19, 2.57154e-19, 
    2.571705e-19, 2.571076e-19, 2.571357e-19, 2.570591e-19, 2.570775e-19, 
    2.570692e-19, 2.570598e-19, 2.570889e-19, 2.57119e-19, 2.571205e-19, 
    2.5713e-19, 2.571554e-19, 2.571103e-19, 2.572564e-19, 2.571646e-19, 
    2.5703e-19, 2.570571e-19, 2.570619e-19, 2.570513e-19, 2.571251e-19, 
    2.570983e-19, 2.571708e-19, 2.571513e-19, 2.571834e-19, 2.571674e-19, 
    2.57165e-19, 2.571447e-19, 2.571318e-19, 2.570993e-19, 2.570732e-19, 
    2.570529e-19, 2.570577e-19, 2.5708e-19, 2.57121e-19, 2.571604e-19, 
    2.571517e-19, 2.57181e-19, 2.571049e-19, 2.571364e-19, 2.571239e-19, 
    2.571565e-19, 2.570861e-19, 2.571435e-19, 2.57071e-19, 2.570776e-19, 
    2.570977e-19, 2.571379e-19, 2.571481e-19, 2.571574e-19, 2.571518e-19, 
    2.571222e-19, 2.571177e-19, 2.570975e-19, 2.570915e-19, 2.570763e-19, 
    2.570633e-19, 2.570749e-19, 2.57087e-19, 2.571226e-19, 2.571542e-19, 
    2.571891e-19, 2.571979e-19, 2.572367e-19, 2.57204e-19, 2.572568e-19, 
    2.572102e-19, 2.572918e-19, 2.571481e-19, 2.572105e-19, 2.57099e-19, 
    2.571111e-19, 2.571323e-19, 2.571827e-19, 2.571564e-19, 2.571876e-19, 
    2.571176e-19, 2.570804e-19, 2.570717e-19, 2.57054e-19, 2.570721e-19, 
    2.570707e-19, 2.570881e-19, 2.570826e-19, 2.571238e-19, 2.571017e-19, 
    2.571647e-19, 2.571876e-19, 2.572532e-19, 2.57293e-19, 2.57335e-19, 
    2.573531e-19, 2.573586e-19, 2.573609e-19 ;

 MEG_acetone =
  8.55093e-17, 8.551773e-17, 8.551619e-17, 8.552264e-17, 8.551913e-17, 
    8.55233e-17, 8.551102e-17, 8.551798e-17, 8.551346e-17, 8.551013e-17, 
    8.553494e-17, 8.552295e-17, 8.554818e-17, 8.554038e-17, 8.556021e-17, 
    8.554687e-17, 8.556293e-17, 8.556e-17, 8.556927e-17, 8.556663e-17, 
    8.557813e-17, 8.55705e-17, 8.558439e-17, 8.55764e-17, 8.557758e-17, 
    8.557022e-17, 8.552553e-17, 8.553339e-17, 8.552502e-17, 8.552615e-17, 
    8.552568e-17, 8.551914e-17, 8.551573e-17, 8.55088e-17, 8.551003e-17, 
    8.551527e-17, 8.552666e-17, 8.552291e-17, 8.553272e-17, 8.553251e-17, 
    8.554332e-17, 8.553844e-17, 8.555679e-17, 8.555162e-17, 8.556674e-17, 
    8.556291e-17, 8.556653e-17, 8.556546e-17, 8.556654e-17, 8.556093e-17, 
    8.556332e-17, 8.555845e-17, 8.553932e-17, 8.554489e-17, 8.552823e-17, 
    8.551797e-17, 8.551128e-17, 8.550663e-17, 8.550729e-17, 8.550851e-17, 
    8.551529e-17, 8.552154e-17, 8.552624e-17, 8.552936e-17, 8.553247e-17, 
    8.554141e-17, 8.554656e-17, 8.555775e-17, 8.555588e-17, 8.555917e-17, 
    8.556253e-17, 8.556798e-17, 8.55671e-17, 8.556947e-17, 8.55592e-17, 
    8.556596e-17, 8.555478e-17, 8.555782e-17, 8.553271e-17, 8.552395e-17, 
    8.551972e-17, 8.551647e-17, 8.550778e-17, 8.551352e-17, 8.551125e-17, 
    8.551711e-17, 8.552056e-17, 8.551887e-17, 8.552945e-17, 8.552531e-17, 
    8.554685e-17, 8.553757e-17, 8.556214e-17, 8.555628e-17, 8.556357e-17, 
    8.555988e-17, 8.556616e-17, 8.556051e-17, 8.557039e-17, 8.557248e-17, 
    8.557104e-17, 8.557677e-17, 8.556017e-17, 8.556647e-17, 8.55188e-17, 
    8.551907e-17, 8.55204e-17, 8.551455e-17, 8.551391e-17, 8.550874e-17, 
    8.551339e-17, 8.551565e-17, 8.55208e-17, 8.552374e-17, 8.552657e-17, 
    8.553281e-17, 8.553969e-17, 8.554951e-17, 8.555665e-17, 8.556142e-17, 
    8.555853e-17, 8.556107e-17, 8.555822e-17, 8.55569e-17, 8.557166e-17, 
    8.556331e-17, 8.557594e-17, 8.557527e-17, 8.55695e-17, 8.557534e-17, 
    8.551927e-17, 8.55177e-17, 8.551173e-17, 8.551647e-17, 8.550818e-17, 
    8.551256e-17, 8.551537e-17, 8.552527e-17, 8.55276e-17, 8.552956e-17, 
    8.553359e-17, 8.553869e-17, 8.554761e-17, 8.555548e-17, 8.556276e-17, 
    8.556223e-17, 8.556241e-17, 8.556397e-17, 8.556002e-17, 8.556463e-17, 
    8.556535e-17, 8.556338e-17, 8.557517e-17, 8.557181e-17, 8.557525e-17, 
    8.557308e-17, 8.551823e-17, 8.55209e-17, 8.551944e-17, 8.552214e-17, 
    8.552019e-17, 8.55287e-17, 8.553126e-17, 8.554338e-17, 8.553855e-17, 
    8.554642e-17, 8.55394e-17, 8.55406e-17, 8.554642e-17, 8.553981e-17, 
    8.555493e-17, 8.554446e-17, 8.556403e-17, 8.555333e-17, 8.556469e-17, 
    8.556272e-17, 8.556604e-17, 8.556896e-17, 8.557275e-17, 8.557956e-17, 
    8.5578e-17, 8.55838e-17, 8.552494e-17, 8.552836e-17, 8.552817e-17, 
    8.553183e-17, 8.553451e-17, 8.554046e-17, 8.55499e-17, 8.55464e-17, 
    8.555297e-17, 8.555425e-17, 8.554433e-17, 8.555031e-17, 8.553073e-17, 
    8.553377e-17, 8.553204e-17, 8.552514e-17, 8.554705e-17, 8.553572e-17, 
    8.555675e-17, 8.555063e-17, 8.556853e-17, 8.555951e-17, 8.557712e-17, 
    8.558437e-17, 8.559174e-17, 8.559975e-17, 8.553034e-17, 8.552801e-17, 
    8.55323e-17, 8.553801e-17, 8.554366e-17, 8.555098e-17, 8.55518e-17, 
    8.555313e-17, 8.555675e-17, 8.555972e-17, 8.555345e-17, 8.556049e-17, 
    8.553425e-17, 8.554808e-17, 8.552702e-17, 8.55332e-17, 8.553773e-17, 
    8.553586e-17, 8.554602e-17, 8.554838e-17, 8.555791e-17, 8.555305e-17, 
    8.558248e-17, 8.556942e-17, 8.560623e-17, 8.559584e-17, 8.552717e-17, 
    8.553039e-17, 8.554145e-17, 8.553621e-17, 8.555153e-17, 8.555526e-17, 
    8.555839e-17, 8.55622e-17, 8.55627e-17, 8.556498e-17, 8.556123e-17, 
    8.556487e-17, 8.5551e-17, 8.555721e-17, 8.554032e-17, 8.554437e-17, 
    8.554255e-17, 8.554047e-17, 8.554688e-17, 8.555352e-17, 8.555384e-17, 
    8.555594e-17, 8.556154e-17, 8.55516e-17, 8.558383e-17, 8.556358e-17, 
    8.55339e-17, 8.553986e-17, 8.554094e-17, 8.553858e-17, 8.555488e-17, 
    8.554895e-17, 8.556495e-17, 8.556066e-17, 8.556773e-17, 8.55642e-17, 
    8.556367e-17, 8.555918e-17, 8.555634e-17, 8.554919e-17, 8.554342e-17, 
    8.553895e-17, 8.554e-17, 8.554493e-17, 8.555397e-17, 8.556266e-17, 
    8.556073e-17, 8.55672e-17, 8.555041e-17, 8.555735e-17, 8.555461e-17, 
    8.55618e-17, 8.554626e-17, 8.555893e-17, 8.554295e-17, 8.55444e-17, 
    8.554883e-17, 8.55577e-17, 8.555994e-17, 8.556199e-17, 8.556076e-17, 
    8.555423e-17, 8.555325e-17, 8.554877e-17, 8.554745e-17, 8.55441e-17, 
    8.554123e-17, 8.55438e-17, 8.554646e-17, 8.555431e-17, 8.556129e-17, 
    8.556898e-17, 8.557093e-17, 8.557947e-17, 8.557226e-17, 8.558391e-17, 
    8.557363e-17, 8.559163e-17, 8.555994e-17, 8.557369e-17, 8.55491e-17, 
    8.555179e-17, 8.555646e-17, 8.556758e-17, 8.556176e-17, 8.556865e-17, 
    8.555322e-17, 8.554501e-17, 8.554309e-17, 8.553918e-17, 8.554319e-17, 
    8.554287e-17, 8.55467e-17, 8.554548e-17, 8.555457e-17, 8.55497e-17, 
    8.556361e-17, 8.556864e-17, 8.558312e-17, 8.559191e-17, 8.560116e-17, 
    8.560515e-17, 8.560639e-17, 8.560689e-17 ;

 MEG_carene_3 =
  3.305452e-17, 3.305785e-17, 3.305724e-17, 3.305979e-17, 3.305841e-17, 
    3.306005e-17, 3.305521e-17, 3.305795e-17, 3.305617e-17, 3.305486e-17, 
    3.306465e-17, 3.305991e-17, 3.306987e-17, 3.306679e-17, 3.307461e-17, 
    3.306935e-17, 3.307569e-17, 3.307454e-17, 3.307819e-17, 3.307715e-17, 
    3.308169e-17, 3.307867e-17, 3.308416e-17, 3.3081e-17, 3.308147e-17, 
    3.307857e-17, 3.306093e-17, 3.306403e-17, 3.306073e-17, 3.306117e-17, 
    3.306099e-17, 3.305841e-17, 3.305706e-17, 3.305433e-17, 3.305482e-17, 
    3.305688e-17, 3.306138e-17, 3.30599e-17, 3.306377e-17, 3.306368e-17, 
    3.306795e-17, 3.306603e-17, 3.307327e-17, 3.307122e-17, 3.307719e-17, 
    3.307568e-17, 3.307711e-17, 3.307669e-17, 3.307712e-17, 3.30749e-17, 
    3.307585e-17, 3.307392e-17, 3.306637e-17, 3.306857e-17, 3.306199e-17, 
    3.305795e-17, 3.305531e-17, 3.305347e-17, 3.305373e-17, 3.305421e-17, 
    3.305689e-17, 3.305936e-17, 3.306121e-17, 3.306245e-17, 3.306367e-17, 
    3.30672e-17, 3.306923e-17, 3.307365e-17, 3.307291e-17, 3.30742e-17, 
    3.307553e-17, 3.307768e-17, 3.307733e-17, 3.307827e-17, 3.307421e-17, 
    3.307688e-17, 3.307247e-17, 3.307367e-17, 3.306377e-17, 3.306031e-17, 
    3.305864e-17, 3.305735e-17, 3.305393e-17, 3.305619e-17, 3.305529e-17, 
    3.305761e-17, 3.305896e-17, 3.30583e-17, 3.306248e-17, 3.306085e-17, 
    3.306935e-17, 3.306568e-17, 3.307538e-17, 3.307307e-17, 3.307594e-17, 
    3.307449e-17, 3.307696e-17, 3.307473e-17, 3.307864e-17, 3.307946e-17, 
    3.307889e-17, 3.308115e-17, 3.307461e-17, 3.307709e-17, 3.305828e-17, 
    3.305838e-17, 3.305891e-17, 3.30566e-17, 3.305634e-17, 3.30543e-17, 
    3.305614e-17, 3.305703e-17, 3.305906e-17, 3.306022e-17, 3.306134e-17, 
    3.30638e-17, 3.306652e-17, 3.307039e-17, 3.307321e-17, 3.307509e-17, 
    3.307396e-17, 3.307496e-17, 3.307383e-17, 3.307331e-17, 3.307913e-17, 
    3.307584e-17, 3.308083e-17, 3.308056e-17, 3.307828e-17, 3.308059e-17, 
    3.305846e-17, 3.305784e-17, 3.305548e-17, 3.305736e-17, 3.305408e-17, 
    3.305581e-17, 3.305692e-17, 3.306083e-17, 3.306174e-17, 3.306252e-17, 
    3.306411e-17, 3.306612e-17, 3.306965e-17, 3.307275e-17, 3.307562e-17, 
    3.307541e-17, 3.307549e-17, 3.30761e-17, 3.307454e-17, 3.307636e-17, 
    3.307664e-17, 3.307587e-17, 3.308052e-17, 3.307919e-17, 3.308055e-17, 
    3.307969e-17, 3.305805e-17, 3.30591e-17, 3.305853e-17, 3.305959e-17, 
    3.305883e-17, 3.306218e-17, 3.306319e-17, 3.306797e-17, 3.306607e-17, 
    3.306917e-17, 3.30664e-17, 3.306688e-17, 3.306918e-17, 3.306657e-17, 
    3.307253e-17, 3.30684e-17, 3.307613e-17, 3.30719e-17, 3.307639e-17, 
    3.307561e-17, 3.307692e-17, 3.307807e-17, 3.307956e-17, 3.308225e-17, 
    3.308164e-17, 3.308393e-17, 3.30607e-17, 3.306205e-17, 3.306197e-17, 
    3.306341e-17, 3.306447e-17, 3.306682e-17, 3.307055e-17, 3.306917e-17, 
    3.307176e-17, 3.307226e-17, 3.306835e-17, 3.307071e-17, 3.306298e-17, 
    3.306418e-17, 3.30635e-17, 3.306078e-17, 3.306942e-17, 3.306495e-17, 
    3.307325e-17, 3.307084e-17, 3.30779e-17, 3.307434e-17, 3.308129e-17, 
    3.308415e-17, 3.308706e-17, 3.309022e-17, 3.306283e-17, 3.306191e-17, 
    3.30636e-17, 3.306586e-17, 3.306809e-17, 3.307098e-17, 3.30713e-17, 
    3.307182e-17, 3.307325e-17, 3.307443e-17, 3.307195e-17, 3.307472e-17, 
    3.306437e-17, 3.306983e-17, 3.306152e-17, 3.306396e-17, 3.306574e-17, 
    3.306501e-17, 3.306902e-17, 3.306995e-17, 3.307371e-17, 3.307179e-17, 
    3.308341e-17, 3.307825e-17, 3.309278e-17, 3.308868e-17, 3.306158e-17, 
    3.306285e-17, 3.306722e-17, 3.306514e-17, 3.307119e-17, 3.307266e-17, 
    3.30739e-17, 3.30754e-17, 3.30756e-17, 3.30765e-17, 3.307502e-17, 
    3.307645e-17, 3.307098e-17, 3.307343e-17, 3.306677e-17, 3.306837e-17, 
    3.306764e-17, 3.306682e-17, 3.306935e-17, 3.307197e-17, 3.30721e-17, 
    3.307293e-17, 3.307514e-17, 3.307122e-17, 3.308394e-17, 3.307595e-17, 
    3.306423e-17, 3.306658e-17, 3.306701e-17, 3.306608e-17, 3.307251e-17, 
    3.307017e-17, 3.307648e-17, 3.307479e-17, 3.307759e-17, 3.307619e-17, 
    3.307598e-17, 3.307421e-17, 3.307309e-17, 3.307027e-17, 3.306799e-17, 
    3.306623e-17, 3.306664e-17, 3.306859e-17, 3.307215e-17, 3.307558e-17, 
    3.307482e-17, 3.307737e-17, 3.307075e-17, 3.307349e-17, 3.30724e-17, 
    3.307524e-17, 3.306911e-17, 3.307411e-17, 3.30678e-17, 3.306837e-17, 
    3.307013e-17, 3.307363e-17, 3.307451e-17, 3.307532e-17, 3.307483e-17, 
    3.307226e-17, 3.307187e-17, 3.30701e-17, 3.306958e-17, 3.306826e-17, 
    3.306712e-17, 3.306814e-17, 3.306919e-17, 3.307229e-17, 3.307504e-17, 
    3.307808e-17, 3.307885e-17, 3.308222e-17, 3.307938e-17, 3.308397e-17, 
    3.307991e-17, 3.308702e-17, 3.307451e-17, 3.307994e-17, 3.307023e-17, 
    3.307129e-17, 3.307314e-17, 3.307752e-17, 3.307523e-17, 3.307795e-17, 
    3.307186e-17, 3.306862e-17, 3.306786e-17, 3.306632e-17, 3.30679e-17, 
    3.306777e-17, 3.306928e-17, 3.30688e-17, 3.307239e-17, 3.307047e-17, 
    3.307596e-17, 3.307795e-17, 3.308366e-17, 3.308713e-17, 3.309078e-17, 
    3.309235e-17, 3.309284e-17, 3.309304e-17 ;

 MEG_ethanol =
  1.71279e-18, 1.713045e-18, 1.712998e-18, 1.713193e-18, 1.713087e-18, 
    1.713213e-18, 1.712842e-18, 1.713052e-18, 1.712916e-18, 1.712816e-18, 
    1.713565e-18, 1.713203e-18, 1.713965e-18, 1.713729e-18, 1.714329e-18, 
    1.713926e-18, 1.714411e-18, 1.714323e-18, 1.714603e-18, 1.714523e-18, 
    1.71487e-18, 1.71464e-18, 1.71506e-18, 1.714818e-18, 1.714854e-18, 
    1.714631e-18, 1.713281e-18, 1.713518e-18, 1.713265e-18, 1.713299e-18, 
    1.713285e-18, 1.713087e-18, 1.712984e-18, 1.712775e-18, 1.712812e-18, 
    1.71297e-18, 1.713315e-18, 1.713201e-18, 1.713498e-18, 1.713491e-18, 
    1.713818e-18, 1.713671e-18, 1.714226e-18, 1.714069e-18, 1.714526e-18, 
    1.71441e-18, 1.71452e-18, 1.714487e-18, 1.71452e-18, 1.714351e-18, 
    1.714423e-18, 1.714276e-18, 1.713697e-18, 1.713866e-18, 1.713362e-18, 
    1.713052e-18, 1.71285e-18, 1.71271e-18, 1.71273e-18, 1.712766e-18, 
    1.712971e-18, 1.71316e-18, 1.713302e-18, 1.713396e-18, 1.71349e-18, 
    1.713761e-18, 1.713916e-18, 1.714255e-18, 1.714198e-18, 1.714297e-18, 
    1.714399e-18, 1.714564e-18, 1.714537e-18, 1.714609e-18, 1.714298e-18, 
    1.714503e-18, 1.714165e-18, 1.714257e-18, 1.713498e-18, 1.713233e-18, 
    1.713105e-18, 1.713007e-18, 1.712744e-18, 1.712918e-18, 1.712849e-18, 
    1.713026e-18, 1.71313e-18, 1.713079e-18, 1.713399e-18, 1.713274e-18, 
    1.713925e-18, 1.713644e-18, 1.714387e-18, 1.71421e-18, 1.71443e-18, 
    1.714319e-18, 1.714509e-18, 1.714338e-18, 1.714637e-18, 1.7147e-18, 
    1.714656e-18, 1.714829e-18, 1.714328e-18, 1.714518e-18, 1.713077e-18, 
    1.713085e-18, 1.713125e-18, 1.712949e-18, 1.71293e-18, 1.712773e-18, 
    1.712914e-18, 1.712982e-18, 1.713138e-18, 1.713226e-18, 1.713312e-18, 
    1.713501e-18, 1.713709e-18, 1.714005e-18, 1.714221e-18, 1.714365e-18, 
    1.714278e-18, 1.714355e-18, 1.714269e-18, 1.714229e-18, 1.714675e-18, 
    1.714423e-18, 1.714804e-18, 1.714784e-18, 1.71461e-18, 1.714786e-18, 
    1.713091e-18, 1.713044e-18, 1.712864e-18, 1.713007e-18, 1.712757e-18, 
    1.712889e-18, 1.712973e-18, 1.713273e-18, 1.713343e-18, 1.713402e-18, 
    1.713524e-18, 1.713678e-18, 1.713948e-18, 1.714186e-18, 1.714406e-18, 
    1.71439e-18, 1.714395e-18, 1.714443e-18, 1.714323e-18, 1.714462e-18, 
    1.714484e-18, 1.714425e-18, 1.714781e-18, 1.714679e-18, 1.714783e-18, 
    1.714718e-18, 1.71306e-18, 1.71314e-18, 1.713097e-18, 1.713178e-18, 
    1.713119e-18, 1.713376e-18, 1.713454e-18, 1.71382e-18, 1.713674e-18, 
    1.713912e-18, 1.7137e-18, 1.713736e-18, 1.713912e-18, 1.713712e-18, 
    1.714169e-18, 1.713853e-18, 1.714444e-18, 1.714121e-18, 1.714464e-18, 
    1.714405e-18, 1.714505e-18, 1.714593e-18, 1.714708e-18, 1.714914e-18, 
    1.714867e-18, 1.715042e-18, 1.713263e-18, 1.713366e-18, 1.71336e-18, 
    1.713471e-18, 1.713552e-18, 1.713732e-18, 1.714017e-18, 1.713911e-18, 
    1.71411e-18, 1.714149e-18, 1.713849e-18, 1.71403e-18, 1.713438e-18, 
    1.71353e-18, 1.713477e-18, 1.713269e-18, 1.713931e-18, 1.713589e-18, 
    1.714224e-18, 1.714039e-18, 1.71458e-18, 1.714308e-18, 1.71484e-18, 
    1.715059e-18, 1.715282e-18, 1.715524e-18, 1.713426e-18, 1.713356e-18, 
    1.713485e-18, 1.713658e-18, 1.713829e-18, 1.71405e-18, 1.714075e-18, 
    1.714115e-18, 1.714224e-18, 1.714314e-18, 1.714125e-18, 1.714337e-18, 
    1.713544e-18, 1.713962e-18, 1.713326e-18, 1.713512e-18, 1.713649e-18, 
    1.713593e-18, 1.7139e-18, 1.713971e-18, 1.714259e-18, 1.714112e-18, 
    1.715002e-18, 1.714607e-18, 1.71572e-18, 1.715406e-18, 1.71333e-18, 
    1.713428e-18, 1.713762e-18, 1.713603e-18, 1.714067e-18, 1.714179e-18, 
    1.714274e-18, 1.714389e-18, 1.714404e-18, 1.714473e-18, 1.71436e-18, 
    1.71447e-18, 1.71405e-18, 1.714238e-18, 1.713728e-18, 1.71385e-18, 
    1.713795e-18, 1.713732e-18, 1.713926e-18, 1.714127e-18, 1.714136e-18, 
    1.7142e-18, 1.714369e-18, 1.714069e-18, 1.715043e-18, 1.714431e-18, 
    1.713533e-18, 1.713714e-18, 1.713746e-18, 1.713675e-18, 1.714168e-18, 
    1.713989e-18, 1.714472e-18, 1.714342e-18, 1.714556e-18, 1.714449e-18, 
    1.714433e-18, 1.714298e-18, 1.714212e-18, 1.713996e-18, 1.713821e-18, 
    1.713686e-18, 1.713718e-18, 1.713867e-18, 1.71414e-18, 1.714403e-18, 
    1.714345e-18, 1.71454e-18, 1.714033e-18, 1.714242e-18, 1.71416e-18, 
    1.714377e-18, 1.713907e-18, 1.71429e-18, 1.713807e-18, 1.713851e-18, 
    1.713985e-18, 1.714253e-18, 1.714321e-18, 1.714383e-18, 1.714345e-18, 
    1.714148e-18, 1.714118e-18, 1.713983e-18, 1.713943e-18, 1.713842e-18, 
    1.713755e-18, 1.713833e-18, 1.713913e-18, 1.71415e-18, 1.714361e-18, 
    1.714594e-18, 1.714653e-18, 1.714911e-18, 1.714693e-18, 1.715045e-18, 
    1.714735e-18, 1.715279e-18, 1.714321e-18, 1.714737e-18, 1.713993e-18, 
    1.714074e-18, 1.714215e-18, 1.714552e-18, 1.714376e-18, 1.714584e-18, 
    1.714118e-18, 1.713869e-18, 1.713812e-18, 1.713693e-18, 1.713814e-18, 
    1.713805e-18, 1.713921e-18, 1.713884e-18, 1.714159e-18, 1.714011e-18, 
    1.714432e-18, 1.714584e-18, 1.715021e-18, 1.715287e-18, 1.715566e-18, 
    1.715687e-18, 1.715724e-18, 1.71574e-18 ;

 MEG_formaldehyde =
  3.425581e-19, 3.426089e-19, 3.425996e-19, 3.426386e-19, 3.426174e-19, 
    3.426426e-19, 3.425685e-19, 3.426105e-19, 3.425832e-19, 3.425631e-19, 
    3.42713e-19, 3.426405e-19, 3.427931e-19, 3.427459e-19, 3.428658e-19, 
    3.427851e-19, 3.428822e-19, 3.428645e-19, 3.429205e-19, 3.429045e-19, 
    3.429741e-19, 3.429279e-19, 3.430119e-19, 3.429636e-19, 3.429707e-19, 
    3.429262e-19, 3.426561e-19, 3.427036e-19, 3.42653e-19, 3.426599e-19, 
    3.42657e-19, 3.426175e-19, 3.425968e-19, 3.425551e-19, 3.425625e-19, 
    3.425941e-19, 3.42663e-19, 3.426403e-19, 3.426996e-19, 3.426983e-19, 
    3.427637e-19, 3.427341e-19, 3.428451e-19, 3.428138e-19, 3.429052e-19, 
    3.428821e-19, 3.429039e-19, 3.428975e-19, 3.429041e-19, 3.428701e-19, 
    3.428846e-19, 3.428551e-19, 3.427395e-19, 3.427732e-19, 3.426724e-19, 
    3.426104e-19, 3.4257e-19, 3.42542e-19, 3.425459e-19, 3.425533e-19, 
    3.425942e-19, 3.42632e-19, 3.426604e-19, 3.426793e-19, 3.426981e-19, 
    3.427521e-19, 3.427832e-19, 3.428509e-19, 3.428396e-19, 3.428595e-19, 
    3.428798e-19, 3.429127e-19, 3.429074e-19, 3.429217e-19, 3.428596e-19, 
    3.429005e-19, 3.428329e-19, 3.428513e-19, 3.426995e-19, 3.426466e-19, 
    3.426209e-19, 3.426013e-19, 3.425489e-19, 3.425836e-19, 3.425698e-19, 
    3.426052e-19, 3.42626e-19, 3.426159e-19, 3.426798e-19, 3.426548e-19, 
    3.42785e-19, 3.427289e-19, 3.428774e-19, 3.42842e-19, 3.428861e-19, 
    3.428638e-19, 3.429017e-19, 3.428676e-19, 3.429273e-19, 3.429399e-19, 
    3.429312e-19, 3.429659e-19, 3.428656e-19, 3.429036e-19, 3.426154e-19, 
    3.42617e-19, 3.426251e-19, 3.425897e-19, 3.425859e-19, 3.425547e-19, 
    3.425828e-19, 3.425964e-19, 3.426275e-19, 3.426452e-19, 3.426624e-19, 
    3.427001e-19, 3.427417e-19, 3.42801e-19, 3.428442e-19, 3.428731e-19, 
    3.428556e-19, 3.42871e-19, 3.428537e-19, 3.428457e-19, 3.429349e-19, 
    3.428845e-19, 3.429609e-19, 3.429568e-19, 3.429219e-19, 3.429573e-19, 
    3.426183e-19, 3.426087e-19, 3.425727e-19, 3.426013e-19, 3.425513e-19, 
    3.425778e-19, 3.425946e-19, 3.426545e-19, 3.426686e-19, 3.426805e-19, 
    3.427048e-19, 3.427356e-19, 3.427896e-19, 3.428372e-19, 3.428811e-19, 
    3.42878e-19, 3.428791e-19, 3.428885e-19, 3.428646e-19, 3.428925e-19, 
    3.428968e-19, 3.428849e-19, 3.429562e-19, 3.429359e-19, 3.429567e-19, 
    3.429435e-19, 3.426119e-19, 3.426281e-19, 3.426193e-19, 3.426356e-19, 
    3.426238e-19, 3.426753e-19, 3.426907e-19, 3.42764e-19, 3.427348e-19, 
    3.427824e-19, 3.427399e-19, 3.427472e-19, 3.427824e-19, 3.427424e-19, 
    3.428338e-19, 3.427706e-19, 3.428889e-19, 3.428241e-19, 3.428929e-19, 
    3.428809e-19, 3.429011e-19, 3.429187e-19, 3.429415e-19, 3.429827e-19, 
    3.429733e-19, 3.430084e-19, 3.426525e-19, 3.426732e-19, 3.42672e-19, 
    3.426942e-19, 3.427104e-19, 3.427464e-19, 3.428035e-19, 3.427822e-19, 
    3.42822e-19, 3.428297e-19, 3.427698e-19, 3.428059e-19, 3.426875e-19, 
    3.427059e-19, 3.426955e-19, 3.426538e-19, 3.427862e-19, 3.427177e-19, 
    3.428448e-19, 3.428079e-19, 3.42916e-19, 3.428615e-19, 3.42968e-19, 
    3.430118e-19, 3.430563e-19, 3.431047e-19, 3.426852e-19, 3.426711e-19, 
    3.42697e-19, 3.427316e-19, 3.427657e-19, 3.4281e-19, 3.428149e-19, 
    3.42823e-19, 3.428448e-19, 3.428628e-19, 3.428249e-19, 3.428674e-19, 
    3.427088e-19, 3.427924e-19, 3.426651e-19, 3.427025e-19, 3.427298e-19, 
    3.427185e-19, 3.4278e-19, 3.427942e-19, 3.428519e-19, 3.428224e-19, 
    3.430004e-19, 3.429214e-19, 3.431439e-19, 3.430811e-19, 3.42666e-19, 
    3.426855e-19, 3.427524e-19, 3.427207e-19, 3.428133e-19, 3.428358e-19, 
    3.428547e-19, 3.428778e-19, 3.428808e-19, 3.428946e-19, 3.428719e-19, 
    3.428939e-19, 3.428101e-19, 3.428476e-19, 3.427455e-19, 3.4277e-19, 
    3.42759e-19, 3.427464e-19, 3.427852e-19, 3.428253e-19, 3.428273e-19, 
    3.4284e-19, 3.428738e-19, 3.428137e-19, 3.430086e-19, 3.428862e-19, 
    3.427067e-19, 3.427428e-19, 3.427492e-19, 3.42735e-19, 3.428335e-19, 
    3.427977e-19, 3.428944e-19, 3.428685e-19, 3.429112e-19, 3.428899e-19, 
    3.428867e-19, 3.428595e-19, 3.428423e-19, 3.427991e-19, 3.427642e-19, 
    3.427372e-19, 3.427436e-19, 3.427734e-19, 3.42828e-19, 3.428806e-19, 
    3.428689e-19, 3.42908e-19, 3.428065e-19, 3.428485e-19, 3.428319e-19, 
    3.428753e-19, 3.427814e-19, 3.42858e-19, 3.427614e-19, 3.427702e-19, 
    3.42797e-19, 3.428506e-19, 3.428641e-19, 3.428765e-19, 3.428691e-19, 
    3.428296e-19, 3.428237e-19, 3.427966e-19, 3.427886e-19, 3.427684e-19, 
    3.42751e-19, 3.427666e-19, 3.427827e-19, 3.428301e-19, 3.428723e-19, 
    3.429187e-19, 3.429306e-19, 3.429822e-19, 3.429386e-19, 3.43009e-19, 
    3.429469e-19, 3.430557e-19, 3.428641e-19, 3.429473e-19, 3.427986e-19, 
    3.428148e-19, 3.428431e-19, 3.429103e-19, 3.428752e-19, 3.429168e-19, 
    3.428235e-19, 3.427739e-19, 3.427623e-19, 3.427387e-19, 3.427628e-19, 
    3.427609e-19, 3.427841e-19, 3.427767e-19, 3.428317e-19, 3.428022e-19, 
    3.428863e-19, 3.429167e-19, 3.430043e-19, 3.430574e-19, 3.431133e-19, 
    3.431374e-19, 3.431449e-19, 3.431479e-19 ;

 MEG_isoprene =
  2.357503e-19, 2.357924e-19, 2.357848e-19, 2.358167e-19, 2.357993e-19, 
    2.3582e-19, 2.357589e-19, 2.357936e-19, 2.35771e-19, 2.357545e-19, 
    2.358776e-19, 2.358182e-19, 2.359432e-19, 2.359045e-19, 2.360027e-19, 
    2.359366e-19, 2.360162e-19, 2.360017e-19, 2.360475e-19, 2.360344e-19, 
    2.360914e-19, 2.360536e-19, 2.361223e-19, 2.360828e-19, 2.360886e-19, 
    2.360522e-19, 2.35831e-19, 2.358699e-19, 2.358285e-19, 2.358341e-19, 
    2.358318e-19, 2.357994e-19, 2.357825e-19, 2.357478e-19, 2.357539e-19, 
    2.357802e-19, 2.358366e-19, 2.358181e-19, 2.358666e-19, 2.358655e-19, 
    2.359191e-19, 2.358949e-19, 2.359858e-19, 2.359601e-19, 2.36035e-19, 
    2.36016e-19, 2.36034e-19, 2.360286e-19, 2.36034e-19, 2.360063e-19, 
    2.360181e-19, 2.35994e-19, 2.358993e-19, 2.359269e-19, 2.358443e-19, 
    2.357936e-19, 2.357601e-19, 2.357371e-19, 2.357404e-19, 2.357464e-19, 
    2.357803e-19, 2.358112e-19, 2.358345e-19, 2.3585e-19, 2.358654e-19, 
    2.359096e-19, 2.359351e-19, 2.359905e-19, 2.359813e-19, 2.359975e-19, 
    2.360142e-19, 2.360411e-19, 2.360368e-19, 2.360485e-19, 2.359977e-19, 
    2.360312e-19, 2.359758e-19, 2.359909e-19, 2.358666e-19, 2.358232e-19, 
    2.358022e-19, 2.357861e-19, 2.357428e-19, 2.357712e-19, 2.357599e-19, 
    2.357893e-19, 2.358064e-19, 2.357981e-19, 2.358504e-19, 2.358299e-19, 
    2.359366e-19, 2.358906e-19, 2.360122e-19, 2.359832e-19, 2.360193e-19, 
    2.36001e-19, 2.360321e-19, 2.360042e-19, 2.360531e-19, 2.360634e-19, 
    2.360563e-19, 2.360846e-19, 2.360025e-19, 2.360337e-19, 2.357977e-19, 
    2.35799e-19, 2.358056e-19, 2.357767e-19, 2.357732e-19, 2.357475e-19, 
    2.357706e-19, 2.357821e-19, 2.358076e-19, 2.358221e-19, 2.358361e-19, 
    2.35867e-19, 2.359011e-19, 2.359497e-19, 2.359851e-19, 2.360087e-19, 
    2.359944e-19, 2.36007e-19, 2.359928e-19, 2.359863e-19, 2.360593e-19, 
    2.36018e-19, 2.360806e-19, 2.360772e-19, 2.360487e-19, 2.360776e-19, 
    2.358e-19, 2.357922e-19, 2.357623e-19, 2.357862e-19, 2.357448e-19, 
    2.357665e-19, 2.357807e-19, 2.358297e-19, 2.358412e-19, 2.35851e-19, 
    2.358709e-19, 2.358961e-19, 2.359403e-19, 2.359793e-19, 2.360153e-19, 
    2.360127e-19, 2.360136e-19, 2.360213e-19, 2.360017e-19, 2.360246e-19, 
    2.360281e-19, 2.360184e-19, 2.360767e-19, 2.360601e-19, 2.360771e-19, 
    2.360664e-19, 2.357948e-19, 2.358081e-19, 2.358009e-19, 2.358143e-19, 
    2.358046e-19, 2.358467e-19, 2.358593e-19, 2.359194e-19, 2.358955e-19, 
    2.359344e-19, 2.358996e-19, 2.359056e-19, 2.359345e-19, 2.359017e-19, 
    2.359766e-19, 2.359247e-19, 2.360216e-19, 2.359686e-19, 2.360249e-19, 
    2.360151e-19, 2.360316e-19, 2.36046e-19, 2.360647e-19, 2.360984e-19, 
    2.360907e-19, 2.361194e-19, 2.358281e-19, 2.35845e-19, 2.358441e-19, 
    2.358622e-19, 2.358754e-19, 2.359049e-19, 2.359517e-19, 2.359343e-19, 
    2.359668e-19, 2.359732e-19, 2.359241e-19, 2.359537e-19, 2.358567e-19, 
    2.358718e-19, 2.358632e-19, 2.358291e-19, 2.359375e-19, 2.358815e-19, 
    2.359856e-19, 2.359553e-19, 2.360439e-19, 2.359992e-19, 2.360864e-19, 
    2.361223e-19, 2.361587e-19, 2.361983e-19, 2.358548e-19, 2.358433e-19, 
    2.358645e-19, 2.358928e-19, 2.359208e-19, 2.35957e-19, 2.359611e-19, 
    2.359677e-19, 2.359855e-19, 2.360003e-19, 2.359692e-19, 2.360041e-19, 
    2.358742e-19, 2.359427e-19, 2.358384e-19, 2.35869e-19, 2.358914e-19, 
    2.358821e-19, 2.359325e-19, 2.359441e-19, 2.359913e-19, 2.359672e-19, 
    2.361129e-19, 2.360483e-19, 2.362304e-19, 2.36179e-19, 2.358391e-19, 
    2.358551e-19, 2.359098e-19, 2.358839e-19, 2.359597e-19, 2.359782e-19, 
    2.359937e-19, 2.360125e-19, 2.36015e-19, 2.360263e-19, 2.360077e-19, 
    2.360258e-19, 2.359571e-19, 2.359878e-19, 2.359042e-19, 2.359243e-19, 
    2.359152e-19, 2.359049e-19, 2.359367e-19, 2.359696e-19, 2.359712e-19, 
    2.359816e-19, 2.360093e-19, 2.359601e-19, 2.361196e-19, 2.360194e-19, 
    2.358724e-19, 2.35902e-19, 2.359073e-19, 2.358956e-19, 2.359763e-19, 
    2.35947e-19, 2.360261e-19, 2.360049e-19, 2.360399e-19, 2.360224e-19, 
    2.360198e-19, 2.359976e-19, 2.359835e-19, 2.359481e-19, 2.359196e-19, 
    2.358974e-19, 2.359026e-19, 2.359271e-19, 2.359718e-19, 2.360148e-19, 
    2.360053e-19, 2.360373e-19, 2.359542e-19, 2.359885e-19, 2.35975e-19, 
    2.360105e-19, 2.359337e-19, 2.359964e-19, 2.359172e-19, 2.359244e-19, 
    2.359464e-19, 2.359903e-19, 2.360013e-19, 2.360115e-19, 2.360054e-19, 
    2.359731e-19, 2.359682e-19, 2.359461e-19, 2.359395e-19, 2.359229e-19, 
    2.359087e-19, 2.359215e-19, 2.359347e-19, 2.359735e-19, 2.36008e-19, 
    2.360461e-19, 2.360557e-19, 2.36098e-19, 2.360624e-19, 2.3612e-19, 
    2.360691e-19, 2.361582e-19, 2.360013e-19, 2.360694e-19, 2.359477e-19, 
    2.35961e-19, 2.359841e-19, 2.360392e-19, 2.360104e-19, 2.360445e-19, 
    2.359681e-19, 2.359274e-19, 2.35918e-19, 2.358986e-19, 2.359184e-19, 
    2.359168e-19, 2.359358e-19, 2.359298e-19, 2.359748e-19, 2.359507e-19, 
    2.360195e-19, 2.360444e-19, 2.361161e-19, 2.361596e-19, 2.362053e-19, 
    2.362251e-19, 2.362312e-19, 2.362337e-19 ;

 MEG_methanol =
  5.873947e-17, 5.874491e-17, 5.874391e-17, 5.87481e-17, 5.874582e-17, 
    5.874852e-17, 5.874058e-17, 5.874508e-17, 5.874217e-17, 5.874001e-17, 
    5.875608e-17, 5.87483e-17, 5.876468e-17, 5.875961e-17, 5.877248e-17, 
    5.876382e-17, 5.877425e-17, 5.877235e-17, 5.877836e-17, 5.877664e-17, 
    5.87841e-17, 5.877916e-17, 5.878816e-17, 5.878298e-17, 5.878375e-17, 
    5.877897e-17, 5.874997e-17, 5.875508e-17, 5.874964e-17, 5.875038e-17, 
    5.875007e-17, 5.874582e-17, 5.874361e-17, 5.873914e-17, 5.873993e-17, 
    5.874332e-17, 5.875071e-17, 5.874827e-17, 5.875464e-17, 5.87545e-17, 
    5.876152e-17, 5.875835e-17, 5.877026e-17, 5.87669e-17, 5.877671e-17, 
    5.877423e-17, 5.877658e-17, 5.877588e-17, 5.877659e-17, 5.877295e-17, 
    5.87745e-17, 5.877133e-17, 5.875892e-17, 5.876253e-17, 5.875172e-17, 
    5.874506e-17, 5.874075e-17, 5.873773e-17, 5.873815e-17, 5.873895e-17, 
    5.874333e-17, 5.874738e-17, 5.875044e-17, 5.875246e-17, 5.875448e-17, 
    5.876028e-17, 5.876362e-17, 5.877088e-17, 5.876967e-17, 5.87718e-17, 
    5.877399e-17, 5.877752e-17, 5.877695e-17, 5.877848e-17, 5.877182e-17, 
    5.877621e-17, 5.876895e-17, 5.877092e-17, 5.875464e-17, 5.874895e-17, 
    5.87462e-17, 5.874409e-17, 5.873848e-17, 5.87422e-17, 5.874072e-17, 
    5.874451e-17, 5.874674e-17, 5.874565e-17, 5.875252e-17, 5.874983e-17, 
    5.876381e-17, 5.875779e-17, 5.877373e-17, 5.876993e-17, 5.877466e-17, 
    5.877226e-17, 5.877634e-17, 5.877267e-17, 5.877908e-17, 5.878044e-17, 
    5.877951e-17, 5.878323e-17, 5.877246e-17, 5.877654e-17, 5.874561e-17, 
    5.874578e-17, 5.874665e-17, 5.874285e-17, 5.874246e-17, 5.87391e-17, 
    5.874212e-17, 5.874356e-17, 5.87469e-17, 5.874881e-17, 5.875065e-17, 
    5.87547e-17, 5.875916e-17, 5.876553e-17, 5.877017e-17, 5.877327e-17, 
    5.877139e-17, 5.877304e-17, 5.877118e-17, 5.877033e-17, 5.87799e-17, 
    5.877449e-17, 5.878269e-17, 5.878225e-17, 5.87785e-17, 5.87823e-17, 
    5.874591e-17, 5.874489e-17, 5.874104e-17, 5.87441e-17, 5.873874e-17, 
    5.874158e-17, 5.874338e-17, 5.874981e-17, 5.875131e-17, 5.875259e-17, 
    5.87552e-17, 5.875851e-17, 5.876431e-17, 5.876941e-17, 5.877413e-17, 
    5.877379e-17, 5.877391e-17, 5.877492e-17, 5.877235e-17, 5.877534e-17, 
    5.877581e-17, 5.877454e-17, 5.878219e-17, 5.878e-17, 5.878224e-17, 
    5.878082e-17, 5.874524e-17, 5.874697e-17, 5.874602e-17, 5.874778e-17, 
    5.874651e-17, 5.875203e-17, 5.875369e-17, 5.876156e-17, 5.875842e-17, 
    5.876353e-17, 5.875897e-17, 5.875975e-17, 5.876353e-17, 5.875924e-17, 
    5.876905e-17, 5.876226e-17, 5.877496e-17, 5.876801e-17, 5.877538e-17, 
    5.877411e-17, 5.877626e-17, 5.877816e-17, 5.878061e-17, 5.878503e-17, 
    5.878402e-17, 5.878779e-17, 5.874959e-17, 5.875181e-17, 5.875169e-17, 
    5.875406e-17, 5.87558e-17, 5.875966e-17, 5.876579e-17, 5.876351e-17, 
    5.876778e-17, 5.876861e-17, 5.876218e-17, 5.876605e-17, 5.875335e-17, 
    5.875532e-17, 5.87542e-17, 5.874972e-17, 5.876394e-17, 5.875659e-17, 
    5.877023e-17, 5.876627e-17, 5.877788e-17, 5.877202e-17, 5.878345e-17, 
    5.878816e-17, 5.879293e-17, 5.879813e-17, 5.87531e-17, 5.875158e-17, 
    5.875436e-17, 5.875807e-17, 5.876174e-17, 5.876649e-17, 5.876702e-17, 
    5.876789e-17, 5.877023e-17, 5.877216e-17, 5.876809e-17, 5.877266e-17, 
    5.875563e-17, 5.876461e-17, 5.875095e-17, 5.875495e-17, 5.875789e-17, 
    5.875668e-17, 5.876327e-17, 5.87648e-17, 5.877099e-17, 5.876783e-17, 
    5.878693e-17, 5.877846e-17, 5.880234e-17, 5.879559e-17, 5.875104e-17, 
    5.875313e-17, 5.876031e-17, 5.87569e-17, 5.876685e-17, 5.876926e-17, 
    5.87713e-17, 5.877377e-17, 5.877409e-17, 5.877557e-17, 5.877314e-17, 
    5.87755e-17, 5.87665e-17, 5.877053e-17, 5.875958e-17, 5.87622e-17, 
    5.876101e-17, 5.875967e-17, 5.876383e-17, 5.876814e-17, 5.876835e-17, 
    5.876971e-17, 5.877334e-17, 5.876689e-17, 5.878781e-17, 5.877467e-17, 
    5.87554e-17, 5.875928e-17, 5.875997e-17, 5.875844e-17, 5.876902e-17, 
    5.876517e-17, 5.877555e-17, 5.877277e-17, 5.877736e-17, 5.877507e-17, 
    5.877472e-17, 5.877181e-17, 5.876996e-17, 5.876533e-17, 5.876158e-17, 
    5.875868e-17, 5.875936e-17, 5.876257e-17, 5.876843e-17, 5.877407e-17, 
    5.877282e-17, 5.877701e-17, 5.876612e-17, 5.877063e-17, 5.876885e-17, 
    5.877351e-17, 5.876343e-17, 5.877165e-17, 5.876128e-17, 5.876222e-17, 
    5.87651e-17, 5.877085e-17, 5.87723e-17, 5.877364e-17, 5.877284e-17, 
    5.87686e-17, 5.876796e-17, 5.876505e-17, 5.876419e-17, 5.876202e-17, 
    5.876016e-17, 5.876183e-17, 5.876356e-17, 5.876865e-17, 5.877318e-17, 
    5.877816e-17, 5.877943e-17, 5.878498e-17, 5.87803e-17, 5.878786e-17, 
    5.878119e-17, 5.879287e-17, 5.87723e-17, 5.878123e-17, 5.876527e-17, 
    5.876701e-17, 5.877004e-17, 5.877726e-17, 5.877349e-17, 5.877796e-17, 
    5.876794e-17, 5.876261e-17, 5.876138e-17, 5.875883e-17, 5.876144e-17, 
    5.876122e-17, 5.876371e-17, 5.876292e-17, 5.876882e-17, 5.876566e-17, 
    5.877468e-17, 5.877795e-17, 5.878735e-17, 5.879305e-17, 5.879905e-17, 
    5.880164e-17, 5.880244e-17, 5.880277e-17 ;

 MEG_pinene_a =
  4.866394e-17, 4.866902e-17, 4.866809e-17, 4.867198e-17, 4.866986e-17, 
    4.867238e-17, 4.866498e-17, 4.866917e-17, 4.866645e-17, 4.866444e-17, 
    4.867939e-17, 4.867216e-17, 4.868738e-17, 4.868267e-17, 4.869463e-17, 
    4.868658e-17, 4.869627e-17, 4.86945e-17, 4.870009e-17, 4.86985e-17, 
    4.870543e-17, 4.870083e-17, 4.87092e-17, 4.870438e-17, 4.87051e-17, 
    4.870066e-17, 4.867372e-17, 4.867846e-17, 4.867341e-17, 4.86741e-17, 
    4.867382e-17, 4.866987e-17, 4.866781e-17, 4.866364e-17, 4.866438e-17, 
    4.866754e-17, 4.86744e-17, 4.867214e-17, 4.867806e-17, 4.867792e-17, 
    4.868445e-17, 4.86815e-17, 4.869257e-17, 4.868945e-17, 4.869856e-17, 
    4.869625e-17, 4.869844e-17, 4.869779e-17, 4.869845e-17, 4.869506e-17, 
    4.869651e-17, 4.869357e-17, 4.868203e-17, 4.868539e-17, 4.867534e-17, 
    4.866916e-17, 4.866513e-17, 4.866233e-17, 4.866273e-17, 4.866346e-17, 
    4.866755e-17, 4.867131e-17, 4.867415e-17, 4.867603e-17, 4.86779e-17, 
    4.868329e-17, 4.86864e-17, 4.869314e-17, 4.869202e-17, 4.8694e-17, 
    4.869603e-17, 4.869931e-17, 4.869878e-17, 4.870021e-17, 4.869402e-17, 
    4.869809e-17, 4.869135e-17, 4.869318e-17, 4.867805e-17, 4.867277e-17, 
    4.867022e-17, 4.866826e-17, 4.866303e-17, 4.866649e-17, 4.866511e-17, 
    4.866865e-17, 4.867072e-17, 4.866971e-17, 4.867609e-17, 4.867359e-17, 
    4.868658e-17, 4.868098e-17, 4.869579e-17, 4.869226e-17, 4.869665e-17, 
    4.869443e-17, 4.869821e-17, 4.869481e-17, 4.870076e-17, 4.870202e-17, 
    4.870116e-17, 4.870461e-17, 4.869461e-17, 4.86984e-17, 4.866967e-17, 
    4.866983e-17, 4.867063e-17, 4.866711e-17, 4.866672e-17, 4.86636e-17, 
    4.866641e-17, 4.866776e-17, 4.867087e-17, 4.867264e-17, 4.867435e-17, 
    4.867811e-17, 4.868226e-17, 4.868818e-17, 4.869248e-17, 4.869536e-17, 
    4.869362e-17, 4.869515e-17, 4.869342e-17, 4.869263e-17, 4.870153e-17, 
    4.86965e-17, 4.870411e-17, 4.87037e-17, 4.870023e-17, 4.870375e-17, 
    4.866995e-17, 4.8669e-17, 4.86654e-17, 4.866826e-17, 4.866327e-17, 
    4.866591e-17, 4.866759e-17, 4.867356e-17, 4.867497e-17, 4.867615e-17, 
    4.867858e-17, 4.868165e-17, 4.868703e-17, 4.869177e-17, 4.869616e-17, 
    4.869584e-17, 4.869595e-17, 4.86969e-17, 4.869451e-17, 4.869729e-17, 
    4.869772e-17, 4.869654e-17, 4.870365e-17, 4.870162e-17, 4.870369e-17, 
    4.870238e-17, 4.866932e-17, 4.867093e-17, 4.867005e-17, 4.867168e-17, 
    4.86705e-17, 4.867563e-17, 4.867717e-17, 4.868448e-17, 4.868157e-17, 
    4.868631e-17, 4.868208e-17, 4.868281e-17, 4.868632e-17, 4.868233e-17, 
    4.869144e-17, 4.868513e-17, 4.869693e-17, 4.869047e-17, 4.869733e-17, 
    4.869614e-17, 4.869814e-17, 4.86999e-17, 4.870218e-17, 4.870629e-17, 
    4.870535e-17, 4.870885e-17, 4.867337e-17, 4.867542e-17, 4.867531e-17, 
    4.867751e-17, 4.867913e-17, 4.868272e-17, 4.868841e-17, 4.86863e-17, 
    4.869026e-17, 4.869103e-17, 4.868505e-17, 4.868866e-17, 4.867686e-17, 
    4.867869e-17, 4.867765e-17, 4.867349e-17, 4.868669e-17, 4.867986e-17, 
    4.869254e-17, 4.868885e-17, 4.869964e-17, 4.86942e-17, 4.870482e-17, 
    4.870919e-17, 4.871364e-17, 4.871846e-17, 4.867662e-17, 4.867521e-17, 
    4.86778e-17, 4.868125e-17, 4.868465e-17, 4.868907e-17, 4.868955e-17, 
    4.869036e-17, 4.869254e-17, 4.869434e-17, 4.869055e-17, 4.869479e-17, 
    4.867898e-17, 4.868731e-17, 4.867462e-17, 4.867834e-17, 4.868107e-17, 
    4.867995e-17, 4.868607e-17, 4.868749e-17, 4.869324e-17, 4.869031e-17, 
    4.870805e-17, 4.870018e-17, 4.872237e-17, 4.87161e-17, 4.867471e-17, 
    4.867665e-17, 4.868332e-17, 4.868016e-17, 4.86894e-17, 4.869164e-17, 
    4.869353e-17, 4.869583e-17, 4.869613e-17, 4.86975e-17, 4.869524e-17, 
    4.869744e-17, 4.868908e-17, 4.869282e-17, 4.868264e-17, 4.868508e-17, 
    4.868398e-17, 4.868273e-17, 4.868659e-17, 4.869059e-17, 4.869079e-17, 
    4.869205e-17, 4.869543e-17, 4.868944e-17, 4.870887e-17, 4.869666e-17, 
    4.867877e-17, 4.868236e-17, 4.868301e-17, 4.868159e-17, 4.869141e-17, 
    4.868784e-17, 4.869748e-17, 4.86949e-17, 4.869916e-17, 4.869703e-17, 
    4.869671e-17, 4.869401e-17, 4.869229e-17, 4.868798e-17, 4.86845e-17, 
    4.868181e-17, 4.868244e-17, 4.868542e-17, 4.869087e-17, 4.869611e-17, 
    4.869494e-17, 4.869884e-17, 4.868872e-17, 4.86929e-17, 4.869125e-17, 
    4.869558e-17, 4.868622e-17, 4.869386e-17, 4.868422e-17, 4.868509e-17, 
    4.868777e-17, 4.869311e-17, 4.869446e-17, 4.86957e-17, 4.869496e-17, 
    4.869102e-17, 4.869043e-17, 4.868773e-17, 4.868693e-17, 4.868492e-17, 
    4.868318e-17, 4.868474e-17, 4.868634e-17, 4.869107e-17, 4.869528e-17, 
    4.869991e-17, 4.870109e-17, 4.870624e-17, 4.87019e-17, 4.870891e-17, 
    4.870272e-17, 4.871357e-17, 4.869446e-17, 4.870276e-17, 4.868793e-17, 
    4.868955e-17, 4.869236e-17, 4.869907e-17, 4.869556e-17, 4.869972e-17, 
    4.869041e-17, 4.868546e-17, 4.868431e-17, 4.868195e-17, 4.868436e-17, 
    4.868417e-17, 4.868648e-17, 4.868575e-17, 4.869123e-17, 4.868829e-17, 
    4.869668e-17, 4.869971e-17, 4.870844e-17, 4.871373e-17, 4.871931e-17, 
    4.872172e-17, 4.872246e-17, 4.872277e-17 ;

 MEG_thujene_a =
  1.227149e-18, 1.227273e-18, 1.22725e-18, 1.227345e-18, 1.227293e-18, 
    1.227354e-18, 1.227174e-18, 1.227276e-18, 1.22721e-18, 1.227162e-18, 
    1.227525e-18, 1.227349e-18, 1.227719e-18, 1.227605e-18, 1.227895e-18, 
    1.2277e-18, 1.227935e-18, 1.227892e-18, 1.228028e-18, 1.227989e-18, 
    1.228158e-18, 1.228046e-18, 1.228249e-18, 1.228132e-18, 1.22815e-18, 
    1.228042e-18, 1.227387e-18, 1.227502e-18, 1.22738e-18, 1.227396e-18, 
    1.227389e-18, 1.227293e-18, 1.227243e-18, 1.227142e-18, 1.22716e-18, 
    1.227237e-18, 1.227404e-18, 1.227349e-18, 1.227492e-18, 1.227489e-18, 
    1.227648e-18, 1.227576e-18, 1.227845e-18, 1.227769e-18, 1.227991e-18, 
    1.227935e-18, 1.227988e-18, 1.227972e-18, 1.227988e-18, 1.227906e-18, 
    1.227941e-18, 1.227869e-18, 1.227589e-18, 1.227671e-18, 1.227427e-18, 
    1.227276e-18, 1.227178e-18, 1.22711e-18, 1.22712e-18, 1.227138e-18, 
    1.227237e-18, 1.227329e-18, 1.227397e-18, 1.227443e-18, 1.227489e-18, 
    1.22762e-18, 1.227695e-18, 1.227859e-18, 1.227832e-18, 1.22788e-18, 
    1.227929e-18, 1.228009e-18, 1.227996e-18, 1.228031e-18, 1.22788e-18, 
    1.227979e-18, 1.227816e-18, 1.22786e-18, 1.227492e-18, 1.227364e-18, 
    1.227302e-18, 1.227254e-18, 1.227127e-18, 1.227211e-18, 1.227178e-18, 
    1.227264e-18, 1.227314e-18, 1.22729e-18, 1.227445e-18, 1.227384e-18, 
    1.2277e-18, 1.227563e-18, 1.227923e-18, 1.227838e-18, 1.227944e-18, 
    1.22789e-18, 1.227982e-18, 1.227899e-18, 1.228044e-18, 1.228075e-18, 
    1.228054e-18, 1.228138e-18, 1.227895e-18, 1.227987e-18, 1.227288e-18, 
    1.227292e-18, 1.227312e-18, 1.227226e-18, 1.227217e-18, 1.227141e-18, 
    1.227209e-18, 1.227242e-18, 1.227318e-18, 1.227361e-18, 1.227402e-18, 
    1.227494e-18, 1.227594e-18, 1.227738e-18, 1.227843e-18, 1.227913e-18, 
    1.227871e-18, 1.227908e-18, 1.227866e-18, 1.227847e-18, 1.228063e-18, 
    1.227941e-18, 1.228126e-18, 1.228116e-18, 1.228031e-18, 1.228117e-18, 
    1.227295e-18, 1.227272e-18, 1.227185e-18, 1.227254e-18, 1.227133e-18, 
    1.227197e-18, 1.227238e-18, 1.227383e-18, 1.227417e-18, 1.227446e-18, 
    1.227505e-18, 1.22758e-18, 1.227711e-18, 1.227826e-18, 1.227932e-18, 
    1.227925e-18, 1.227927e-18, 1.22795e-18, 1.227892e-18, 1.22796e-18, 
    1.22797e-18, 1.227942e-18, 1.228114e-18, 1.228065e-18, 1.228115e-18, 
    1.228084e-18, 1.22728e-18, 1.227319e-18, 1.227298e-18, 1.227337e-18, 
    1.227309e-18, 1.227433e-18, 1.227471e-18, 1.227649e-18, 1.227578e-18, 
    1.227693e-18, 1.22759e-18, 1.227608e-18, 1.227693e-18, 1.227596e-18, 
    1.227818e-18, 1.227664e-18, 1.227951e-18, 1.227794e-18, 1.227961e-18, 
    1.227932e-18, 1.227981e-18, 1.228023e-18, 1.228079e-18, 1.228179e-18, 
    1.228156e-18, 1.228241e-18, 1.227378e-18, 1.227428e-18, 1.227426e-18, 
    1.227479e-18, 1.227519e-18, 1.227606e-18, 1.227744e-18, 1.227693e-18, 
    1.227789e-18, 1.227808e-18, 1.227662e-18, 1.22775e-18, 1.227463e-18, 
    1.227508e-18, 1.227482e-18, 1.227381e-18, 1.227702e-18, 1.227536e-18, 
    1.227844e-18, 1.227755e-18, 1.228017e-18, 1.227885e-18, 1.228143e-18, 
    1.228249e-18, 1.228357e-18, 1.228474e-18, 1.227458e-18, 1.227423e-18, 
    1.227486e-18, 1.22757e-18, 1.227653e-18, 1.22776e-18, 1.227772e-18, 
    1.227791e-18, 1.227844e-18, 1.227888e-18, 1.227796e-18, 1.227899e-18, 
    1.227515e-18, 1.227717e-18, 1.227409e-18, 1.227499e-18, 1.227566e-18, 
    1.227538e-18, 1.227687e-18, 1.227722e-18, 1.227862e-18, 1.22779e-18, 
    1.228221e-18, 1.22803e-18, 1.228569e-18, 1.228417e-18, 1.227411e-18, 
    1.227458e-18, 1.22762e-18, 1.227543e-18, 1.227768e-18, 1.227823e-18, 
    1.227868e-18, 1.227924e-18, 1.227932e-18, 1.227965e-18, 1.22791e-18, 
    1.227963e-18, 1.22776e-18, 1.227851e-18, 1.227604e-18, 1.227663e-18, 
    1.227636e-18, 1.227606e-18, 1.2277e-18, 1.227797e-18, 1.227802e-18, 
    1.227833e-18, 1.227915e-18, 1.227769e-18, 1.228241e-18, 1.227945e-18, 
    1.22751e-18, 1.227597e-18, 1.227613e-18, 1.227578e-18, 1.227817e-18, 
    1.22773e-18, 1.227965e-18, 1.227902e-18, 1.228005e-18, 1.227954e-18, 
    1.227946e-18, 1.22788e-18, 1.227838e-18, 1.227734e-18, 1.227649e-18, 
    1.227584e-18, 1.227599e-18, 1.227671e-18, 1.227804e-18, 1.227931e-18, 
    1.227903e-18, 1.227997e-18, 1.227752e-18, 1.227853e-18, 1.227813e-18, 
    1.227918e-18, 1.227691e-18, 1.227876e-18, 1.227642e-18, 1.227663e-18, 
    1.227728e-18, 1.227858e-18, 1.227891e-18, 1.227921e-18, 1.227903e-18, 
    1.227808e-18, 1.227793e-18, 1.227728e-18, 1.227708e-18, 1.227659e-18, 
    1.227617e-18, 1.227655e-18, 1.227694e-18, 1.227809e-18, 1.227911e-18, 
    1.228024e-18, 1.228052e-18, 1.228177e-18, 1.228072e-18, 1.228242e-18, 
    1.228092e-18, 1.228355e-18, 1.227891e-18, 1.228093e-18, 1.227732e-18, 
    1.227772e-18, 1.22784e-18, 1.228003e-18, 1.227918e-18, 1.228019e-18, 
    1.227793e-18, 1.227672e-18, 1.227644e-18, 1.227587e-18, 1.227646e-18, 
    1.227641e-18, 1.227697e-18, 1.227679e-18, 1.227813e-18, 1.227741e-18, 
    1.227945e-18, 1.228019e-18, 1.228231e-18, 1.22836e-18, 1.228495e-18, 
    1.228554e-18, 1.228572e-18, 1.228579e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -4.642471e-25, 4.395241e-25, -1.18122e-25, -5.494041e-26, 1.565805e-25, 
    -5.796222e-25, -4.093066e-25, -2.472314e-26, -4.148007e-25, 
    -2.884375e-25, 2.747026e-25, -1.922916e-25, 5.76876e-26, -3.873304e-25, 
    -5.60393e-25, -1.922916e-25, -1.813036e-25, -5.081995e-25, -9.065174e-26, 
    1.318573e-25, -2.197612e-26, 4.202949e-25, -4.807293e-25, -3.845826e-26, 
    -2.582203e-25, 8.241083e-26, -4.202947e-25, -6.867554e-26, -3.076667e-25, 
    -1.20869e-25, -8.790471e-26, -1.648214e-25, 2.280031e-25, -2.225089e-25, 
    -8.790471e-26, 2.11521e-25, -6.510448e-25, -4.862233e-25, 2.032799e-25, 
    -1.867976e-25, 2.939317e-25, 1.373513e-25, -2.637143e-25, 3.351371e-25, 
    -1.318571e-25, 4.395241e-25, -5.219339e-26, -1.20869e-25, -2.115208e-25, 
    -2.225089e-25, 8.241157e-27, -1.867976e-25, 5.494058e-26, 2.747033e-26, 
    -2.472314e-26, 2.280031e-25, -2.856905e-25, 1.620745e-25, -5.768744e-26, 
    -8.735538e-25, -3.104137e-25, -1.730625e-25, 6.043463e-26, 1.181221e-25, 
    -1.126279e-25, 4.010657e-25, 2.582204e-25, 1.263632e-25, 1.400983e-25, 
    -2.966786e-25, -2.664613e-25, 3.076668e-25, -1.730625e-25, 4.944653e-26, 
    7.169735e-25, -5.851162e-25, -2.032798e-25, 1.922926e-26, 4.120545e-26, 
    3.571133e-25, -2.747024e-25, -9.889281e-26, -1.098809e-25, 2.14268e-25, 
    -3.021719e-26, 7.416975e-26, -2.25256e-25, 3.598603e-25, -4.779822e-25, 
    -1.18122e-25, 5.494132e-27, 5.219355e-26, 1.098818e-26, -1.538333e-25, 
    3.021735e-26, -8.790471e-26, 1.867978e-25, -1.071339e-25, 7.416975e-26, 
    -8.240992e-27, -1.565803e-25, 1.510864e-25, 7.691677e-26, -6.78515e-25, 
    -1.648207e-26, -2.747016e-26, -2.966786e-25, -1.922909e-26, 
    -3.845826e-26, 7.416975e-26, -2.637143e-25, 1.373521e-26, 2.747033e-26, 
    3.543663e-25, -4.697411e-25, 5.494132e-27, -3.46125e-25, -2.389911e-25, 
    2.005329e-25, 1.291103e-25, -1.565803e-25, 2.197628e-26, -1.813036e-25, 
    -2.499792e-25, 1.950388e-25, -6.318156e-25, -4.202947e-25, -4.038125e-25, 
    -1.318571e-25, -3.296421e-26, -2.774494e-25, -1.867976e-25, 
    -5.466578e-25, -1.620744e-25, -2.527262e-25, 4.505122e-25, 1.593275e-25, 
    -2.197619e-25, -3.983185e-25, -2.417381e-25, -2.115208e-25, 2.08774e-25, 
    -2.032798e-25, -4.367769e-25, -2.115208e-25, -4.148007e-25, 
    -9.614578e-26, -8.515768e-26, -5.521519e-25, 2.472331e-26, -6.70274e-25, 
    -5.768744e-26, -2.582203e-25, -2.472321e-25, 1.291103e-25, 6.592867e-26, 
    7.96638e-26, 4.889705e-25, 5.274289e-25, -3.900774e-25, -5.494041e-26, 
    2.362442e-25, -1.593274e-25, -6.565389e-25, -1.098809e-25, -3.296429e-25, 
    2.801966e-25, -2.197612e-26, -8.515768e-26, -2.554732e-25, -9.339876e-26, 
    -1.15375e-25, -5.576459e-25, -2.197612e-26, -3.351369e-25, -4.202947e-25, 
    -6.592851e-26, 3.18655e-25, -4.395231e-26, -2.087738e-25, 5.76876e-26, 
    -4.724882e-25, -3.296421e-26, 1.977859e-25, -6.675269e-25, 3.488722e-25, 
    -1.675684e-25, -4.285358e-25, -4.010655e-25, 1.04387e-25, 3.955716e-25, 
    -6.318148e-26, -4.944636e-26, -5.6314e-25, 2.197628e-26, -5.494041e-26, 
    -3.598602e-25, 2.362442e-25, 4.120538e-25, -2.801964e-25, -4.944636e-26, 
    -3.873304e-25, 4.395248e-26, 2.14268e-25, 1.730626e-25, 3.323901e-25, 
    -2.087738e-25, 1.703156e-25, 3.378841e-25, -3.488721e-25, -1.895446e-25, 
    6.043463e-26, -2.417381e-25, -1.428452e-25, 1.208692e-25, -3.681012e-25, 
    -1.373504e-26, 2.252561e-25, 1.648223e-26, -4.752352e-25, 1.703156e-25, 
    2.719555e-25, 4.944653e-26, 3.763425e-25, -2.747024e-25, -2.829435e-25, 
    -2.911845e-25, -3.845834e-25, 1.181221e-25, 2.08774e-25, -3.351369e-25, 
    -1.922909e-26, 3.571133e-25, -4.395231e-26, -1.950387e-25, 6.043463e-26, 
    -1.373512e-25, -3.104137e-25, -7.966364e-26, 1.922918e-25, -1.675684e-25, 
    -2.829435e-25, -1.675684e-25, 1.922926e-26, -2.197612e-26, -4.395239e-25, 
    1.318573e-25, 1.428454e-25, 2.747107e-27, -2.170149e-25, 2.472331e-26, 
    6.86757e-26, 4.395248e-26, 6.043463e-26, -1.703155e-25, -3.296421e-26, 
    1.208692e-25, 3.845843e-26, -3.241488e-25, -3.516191e-25, -3.076667e-25, 
    -2.554732e-25, 2.08774e-25, 3.571133e-25, 8.790487e-26, -3.131607e-25, 
    -2.884375e-25, 1.922918e-25, 3.159079e-25, -1.922916e-25, 8.790487e-26, 
    -2.856905e-25, -1.840506e-25, -3.186548e-25, 8.241083e-26, -1.483393e-25, 
    -3.296429e-25, 2.197628e-26, 3.26896e-25, -1.867976e-25, -1.098809e-25, 
    -3.186548e-25, -3.214018e-25, -1.15375e-25, 3.351371e-25, -1.400982e-25, 
    8.790487e-26, -1.428452e-25, -2.747024e-25, -6.043446e-26, -8.790471e-26, 
    -1.071339e-25, 8.515785e-26, -3.214018e-25, -6.318148e-26, -6.345626e-25, 
    1.098818e-26, 2.08774e-25, 2.225091e-25, -7.691661e-26, 2.856907e-25, 
    -6.318148e-26, 1.428454e-25, 1.510864e-25, 3.296438e-26, 4.944653e-26, 
    7.96638e-26, -7.142256e-26, 3.159079e-25, 3.021728e-25, -3.43378e-25, 
    -3.076667e-25, -1.15375e-25, 9.339892e-26, -3.845826e-26, 1.263632e-25, 
    2.609674e-25, -1.18122e-25, -1.813036e-25, -1.016398e-25, 4.257889e-25, 
    -3.845826e-26, 2.856907e-25, 1.428454e-25, 2.08774e-25, -2.225089e-25, 
    1.373521e-26, -2.36244e-25, 1.922918e-25, 6.86757e-26, 1.510864e-25, 
    -5.60393e-25, 1.922918e-25, -3.983185e-25, 3.735955e-25, -5.246816e-25, 
    6.977444e-25, -5.493967e-27 ;

 M_LITR2C_TO_LEACHING =
  -3.021727e-25, -1.043869e-25, -1.18122e-25, 9.065187e-26, -1.291101e-25, 
    2.087739e-25, -2.554732e-25, 1.510864e-25, 1.126281e-25, 9.889295e-26, 
    -7.691664e-26, -3.845829e-26, 2.087739e-25, 1.703156e-25, -2.801965e-25, 
    5.351392e-32, 2.582204e-25, -6.592854e-26, -1.098809e-25, 1.455924e-25, 
    -1.922917e-25, -2.197614e-26, 1.64822e-26, 2.801966e-25, 2.197625e-26, 
    1.153751e-25, -6.592854e-26, 5.494055e-26, -2.911846e-25, 1.208691e-25, 
    1.64822e-26, -2.197614e-26, 6.867567e-26, -1.813036e-25, -1.620744e-25, 
    6.04346e-26, 5.351406e-32, 1.04387e-25, 3.955716e-25, 1.04387e-25, 
    -7.142259e-26, 2.362442e-25, -5.493996e-27, -6.592854e-26, 2.197625e-26, 
    -3.845829e-26, -2.527262e-25, 3.84584e-26, -2.692084e-25, -1.043869e-25, 
    1.64822e-26, 1.922918e-25, -2.197614e-26, -4.944639e-26, -8.790474e-26, 
    6.592865e-26, -8.241021e-27, 1.538334e-25, 8.241128e-27, -1.016399e-25, 
    -1.098805e-26, 3.84584e-26, 8.515782e-26, -5.494044e-26, 2.17015e-25, 
    -9.889284e-26, -1.648209e-26, 2.14268e-25, -5.493996e-27, 6.015985e-25, 
    -3.296429e-25, 1.730626e-25, 7.691675e-26, -7.966367e-26, -2.389911e-25, 
    8.24108e-26, -1.648209e-26, 5.494103e-27, -8.241069e-26, 2.692085e-25, 
    1.318572e-25, 3.84584e-26, -3.296424e-26, 1.510864e-25, 2.472323e-25, 
    1.04387e-25, 1.126281e-25, -2.499792e-25, -5.768747e-26, 1.09881e-25, 
    5.351392e-32, 2.856906e-25, -2.197614e-26, 5.351386e-32, 4.94465e-26, 
    -2.197619e-25, -9.614581e-26, 3.84584e-26, 1.455924e-25, -2.197619e-25, 
    -1.043869e-25, -2.527262e-25, 1.098815e-26, 8.24108e-26, -7.691664e-26, 
    -1.098805e-26, -9.339879e-26, 1.0164e-25, -2.856905e-25, 5.351417e-32, 
    5.494103e-27, 8.24108e-26, -2.197619e-25, -3.845829e-26, -2.444852e-25, 
    -1.840506e-25, 1.703156e-25, 8.790485e-26, 9.339889e-26, 2.087739e-25, 
    -2.28003e-25, -4.944639e-26, 1.483394e-25, -1.648209e-26, 1.07134e-25, 
    -7.966367e-26, 1.04387e-25, -6.318152e-26, 2.417382e-25, 1.703156e-25, 
    7.14227e-26, 5.219352e-26, 5.494055e-26, -6.867557e-26, 6.592865e-26, 
    1.703156e-25, -4.395234e-26, -4.395234e-26, -1.400982e-25, 5.351403e-32, 
    7.14227e-26, 4.669947e-26, -3.900775e-25, 1.758096e-25, -3.021722e-26, 
    -1.12628e-25, 5.351382e-32, 9.339889e-26, -2.389911e-25, 1.181221e-25, 
    -5.494044e-26, -2.74702e-26, -1.813036e-25, -9.614581e-26, -2.444852e-25, 
    -8.241021e-27, 1.483394e-25, 2.19762e-25, -3.928245e-25, 1.263632e-25, 
    -1.263631e-25, -8.790474e-26, 1.318572e-25, 2.19762e-25, 7.14227e-26, 
    7.691675e-26, -1.867976e-25, -3.186548e-25, -1.455923e-25, 8.24108e-26, 
    1.153751e-25, 1.09881e-25, 8.24108e-26, -2.444852e-25, -1.428452e-25, 
    3.21402e-25, -2.692084e-25, 5.768757e-26, 1.867977e-25, 5.351371e-32, 
    1.318572e-25, 1.840507e-25, 1.04387e-25, -2.060268e-25, -4.175477e-25, 
    -4.944639e-26, -2.582203e-25, -3.021722e-26, -4.944639e-26, 5.494055e-26, 
    2.087739e-25, -1.977857e-25, 4.120543e-26, 1.263632e-25, -2.417381e-25, 
    6.04346e-26, 2.966787e-25, -3.186548e-25, -1.977857e-25, 1.813037e-25, 
    -8.241021e-27, 7.691675e-26, 4.395245e-26, 9.889295e-26, 1.64822e-26, 
    -2.25256e-25, -1.098805e-26, -7.691664e-26, 7.14227e-26, 4.42271e-25, 
    -2.582203e-25, 7.14227e-26, 2.74703e-26, 2.197625e-26, 2.14268e-25, 
    1.703156e-25, 1.922923e-26, 9.339889e-26, -9.889284e-26, -1.538333e-25, 
    -6.592854e-26, 1.346043e-25, 1.483394e-25, 5.219352e-26, -9.065177e-26, 
    -1.373512e-25, -6.592854e-26, -3.571132e-25, -3.681013e-25, 1.373518e-26, 
    5.494103e-27, 8.24108e-26, -6.592854e-26, 1.648215e-25, 5.494103e-27, 
    1.153751e-25, 2.747078e-27, -1.20869e-25, 1.64822e-26, -2.28003e-25, 
    6.04346e-26, -2.197619e-25, -2.801965e-25, -3.845829e-26, -1.950387e-25, 
    -2.362441e-25, 4.94465e-26, -1.373507e-26, 7.691675e-26, -1.867976e-25, 
    -1.373512e-25, -4.395234e-26, -2.032798e-25, 1.64822e-26, 1.04387e-25, 
    -1.648214e-25, 7.966377e-26, 6.04346e-26, -2.74702e-26, 5.219352e-26, 
    -2.499792e-25, -1.758095e-25, -2.472317e-26, 2.472328e-26, 2.19762e-25, 
    -3.571127e-26, -2.472317e-26, 3.26896e-25, -2.142679e-25, -1.428452e-25, 
    1.04387e-25, -9.339879e-26, -5.493996e-27, 7.966377e-26, 1.236162e-25, 
    -4.395234e-26, -1.593274e-25, 2.527263e-25, 1.840507e-25, -8.241021e-27, 
    -1.977857e-25, -7.691664e-26, 1.593275e-25, 1.236162e-25, -3.983186e-25, 
    -1.538333e-25, 3.104139e-25, 1.236162e-25, 1.538334e-25, -1.922917e-25, 
    1.64822e-26, 2.966787e-25, 5.494103e-27, 1.318572e-25, -9.065177e-26, 
    9.889295e-26, 1.730626e-25, -2.499792e-25, 2.197625e-26, -7.416961e-26, 
    1.730626e-25, -1.675685e-25, -7.691664e-26, 9.889295e-26, -9.889284e-26, 
    3.571138e-26, -2.115208e-25, 2.087739e-25, -5.494044e-26, 1.400983e-25, 
    -2.142679e-25, -9.339879e-26, 2.74703e-26, -1.785566e-25, -2.197614e-26, 
    -2.719554e-25, -8.515771e-26, 9.889295e-26, -1.922917e-25, -2.637143e-25, 
    -1.373512e-25, 3.296435e-26, 4.94465e-26, 1.813037e-25, 2.17015e-25, 
    -6.592854e-26, -2.197614e-26, 8.790485e-26, -1.263631e-25, 9.339889e-26, 
    -3.296424e-26, 1.153751e-25, -2.74702e-26, -3.021722e-26, 2.14268e-25, 
    -4.395234e-26, 6.867567e-26, -3.021727e-25 ;

 M_LITR3C_TO_LEACHING =
  -1.043869e-25, -3.159076e-26, -2.747022e-26, 5.494052e-26, -1.922917e-25, 
    -6.592857e-26, 5.494076e-27, -3.57113e-26, -1.263631e-25, 3.983189e-26, 
    -1.071339e-25, 1.098813e-26, -3.708481e-26, -1.098807e-26, -2.747022e-26, 
    2.060271e-26, -1.37351e-26, -1.09881e-25, -9.065179e-26, -6.730208e-26, 
    1.524599e-25, -5.219344e-26, -1.332307e-25, 4.944647e-26, -5.494047e-26, 
    -1.510863e-25, -1.648215e-25, -5.768749e-26, 8.790482e-26, -5.081993e-26, 
    2.197622e-26, 3.296432e-26, -2.170149e-25, 3.296432e-26, -2.28003e-25, 
    -5.494023e-27, -3.296427e-26, 1.304837e-25, -7.829018e-26, -2.334968e-26, 
    1.030135e-25, -5.494047e-26, -8.241047e-27, -3.983183e-26, 1.263632e-25, 
    -2.747022e-26, -8.653126e-26, 1.510866e-26, -3.021725e-26, -5.768749e-26, 
    -9.20253e-26, -1.236158e-26, -8.241071e-26, 8.378428e-26, -8.790477e-26, 
    -1.12628e-25, 8.790482e-26, -8.515774e-26, 6.180808e-26, -1.277366e-25, 
    -1.15375e-25, -8.10372e-26, 2.197622e-26, 1.744361e-25, -1.194956e-25, 
    1.373515e-26, 8.378428e-26, -6.592857e-26, -1.922915e-26, -2.47232e-26, 
    1.09881e-25, -1.016399e-25, -6.592857e-26, 8.790482e-26, -5.356696e-26, 
    4.669945e-26, 2.747028e-26, 1.07134e-25, -6.867559e-26, 4.807296e-26, 
    -2.197617e-26, 1.840507e-25, -4.669939e-26, -9.61456e-27, -1.263631e-25, 
    1.09881e-25, -1.400982e-25, -3.57113e-26, 7.691672e-26, -9.339881e-26, 
    1.730626e-25, 1.016399e-25, 7.691672e-26, 5.494076e-27, -6.455506e-26, 
    5.356701e-26, -1.098807e-26, -3.296427e-26, 1.565804e-25, -7.142262e-26, 
    1.098813e-26, -2.197617e-26, 6.31816e-26, -8.241047e-27, 8.241101e-27, 
    2.472325e-26, -8.241071e-26, -1.12628e-25, -4.807291e-26, -9.477233e-26, 
    2.747052e-27, 1.510864e-25, -1.428453e-25, 4.807296e-26, -4.807291e-26, 
    -1.304836e-25, -1.236158e-26, -2.746998e-27, 3.159081e-26, -5.768749e-26, 
    -9.751935e-26, -3.021725e-26, 1.950388e-25, 9.614614e-27, 8.790482e-26, 
    1.400983e-25, -7.142262e-26, -4.944642e-26, 3.708486e-26, 7.416969e-26, 
    -3.845832e-26, -2.747022e-26, 5.494052e-26, -1.236158e-26, 1.455923e-25, 
    -9.614584e-26, -1.400982e-25, -1.291101e-25, -7.966369e-26, 7.416969e-26, 
    1.167486e-25, 5.21935e-26, 3.845837e-26, 2.747028e-26, -7.279613e-26, 
    -2.060266e-26, 2.747028e-26, -1.648215e-25, 4.120564e-27, -6.867559e-26, 
    -7.142262e-26, 7.142267e-26, -6.867559e-26, 5.21935e-26, 9.065185e-26, 
    -1.373512e-25, -1.071339e-25, -5.494047e-26, 4.395242e-26, -2.197617e-26, 
    -1.12628e-25, 8.103726e-26, -8.241047e-27, -6.043452e-26, 8.378428e-26, 
    1.92292e-26, -1.236161e-25, -1.09881e-25, -9.889287e-26, -1.016399e-25, 
    -8.241047e-27, -4.807291e-26, 4.669945e-26, -1.922915e-26, 1.098813e-26, 
    -1.922915e-26, -1.318572e-25, 1.648217e-26, -3.845832e-26, -9.614584e-26, 
    1.840507e-25, -2.499792e-25, 2.747028e-26, -2.747022e-26, 2.472325e-26, 
    -1.867977e-25, 8.378428e-26, 2.472325e-26, 4.807296e-26, 4.807296e-26, 
    6.867589e-27, 2.675693e-32, -8.927828e-26, 3.708486e-26, 3.983189e-26, 
    -1.607009e-25, -7.279613e-26, -1.346042e-25, 1.455923e-25, 1.455923e-25, 
    8.241101e-27, 8.241101e-27, 1.04387e-25, -5.631398e-26, 3.571135e-26, 
    -1.18122e-25, -4.395237e-26, 8.241101e-27, -5.768749e-26, 1.236164e-26, 
    -1.071339e-25, -8.10372e-26, 4.669945e-26, 2.747052e-27, 1.92292e-26, 
    -8.241047e-27, 9.614589e-26, 3.983189e-26, -1.37351e-26, -1.675685e-25, 
    -5.356696e-26, -7.829018e-26, -1.785566e-25, 1.854242e-25, -2.746998e-27, 
    -4.944642e-26, -5.768749e-26, 2.675695e-32, -6.592857e-26, -9.065179e-26, 
    3.02173e-26, 3.296432e-26, -1.675685e-25, 3.433784e-26, -7.554316e-26, 
    -4.944642e-26, 1.785566e-25, -5.768749e-26, 4.395242e-26, -1.620744e-25, 
    2.675692e-32, 5.631404e-26, -2.197617e-26, -4.257886e-26, -1.208691e-25, 
    -1.648212e-26, -8.515774e-26, 3.296432e-26, 1.57954e-25, 1.346042e-25, 
    -1.37351e-26, -4.395237e-26, 1.428453e-25, 8.653131e-26, -8.10372e-26, 
    -5.631398e-26, -3.296427e-26, -6.730208e-26, -2.884373e-26, 
    -1.373486e-27, -6.592857e-26, 4.12054e-26, -7.142262e-26, 8.103726e-26, 
    -1.09881e-25, 9.477238e-26, -2.087739e-25, 1.373515e-26, 9.614589e-26, 
    -7.691667e-26, -8.241047e-27, -7.142262e-26, 1.153751e-25, -7.416964e-26, 
    -1.15375e-25, -1.400982e-25, -2.156414e-25, -9.20253e-26, -7.691667e-26, 
    -7.829018e-26, 5.494076e-27, 1.098813e-26, -6.592857e-26, -1.222426e-25, 
    -9.339881e-26, 6.867565e-26, -1.37351e-26, -3.845832e-26, 9.202536e-26, 
    2.747052e-27, -1.18122e-25, -2.746998e-27, 1.373515e-26, -1.291101e-25, 
    -5.219344e-26, -8.927828e-26, -6.318154e-26, 4.12054e-26, 3.571135e-26, 
    2.747028e-26, 8.515779e-26, -6.867559e-26, -5.906101e-26, -3.57113e-26, 
    -4.120535e-26, 1.016399e-25, 2.675688e-32, -6.043452e-26, -9.477233e-26, 
    3.296432e-26, 6.730214e-26, -4.120535e-26, 1.167486e-25, -8.790477e-26, 
    2.472325e-26, -4.120535e-26, 1.675685e-25, 6.043457e-26, -2.197617e-26, 
    -3.021725e-26, 3.02173e-26, -2.746998e-27, -6.867559e-26, -1.263631e-25, 
    -4.944642e-26, -5.494047e-26, -1.167485e-25, -1.140015e-25, 
    -1.648212e-26, 3.02173e-26, 1.291102e-25, 3.845837e-26, -1.236158e-26, 
    -6.318154e-26, -7.279613e-26, -2.060266e-26, -7.554316e-26, -1.016399e-25 ;

 M_SOIL1C_TO_LEACHING =
  -2.208014e-20, -3.02242e-20, 2.566799e-20, 1.942908e-21, 5.434642e-21, 
    -1.145039e-22, 1.698563e-20, -2.067601e-21, -1.905096e-20, -1.189759e-20, 
    -1.626435e-20, 1.4507e-21, -2.053673e-20, 2.278527e-20, 1.458296e-20, 
    4.508733e-20, -5.297531e-21, 4.957995e-20, -1.328015e-20, -1.256231e-20, 
    1.767294e-20, 2.470389e-20, 1.525247e-20, -2.605139e-20, 2.148189e-20, 
    -1.838032e-20, 4.159223e-20, -4.119274e-20, 3.133702e-20, -1.660363e-20, 
    1.744434e-21, 2.298049e-21, 4.871029e-20, -3.996116e-21, 2.076713e-20, 
    -1.494033e-20, -3.470717e-20, 1.202254e-20, -8.761833e-21, 3.596167e-20, 
    -2.480569e-20, 1.13655e-20, -3.905898e-20, -9.158504e-21, -3.381657e-20, 
    2.643268e-21, 3.586158e-20, 1.795764e-20, 1.120036e-20, 1.640716e-20, 
    -1.204377e-20, 6.850511e-22, -1.544301e-20, 7.953217e-21, -8.555726e-21, 
    -2.293936e-20, 4.066942e-20, -4.970689e-21, -1.902186e-20, 3.164859e-20, 
    4.188288e-20, 3.319711e-20, -3.010685e-20, 3.582991e-20, 7.388018e-21, 
    -1.422843e-20, -3.913418e-20, -2.730672e-20, -1.886324e-20, 
    -7.615918e-20, 1.910667e-21, -2.918544e-20, 3.211481e-20, -3.33775e-20, 
    2.067949e-20, -1.432881e-20, -3.048403e-20, 2.128696e-21, -7.360617e-21, 
    -2.60309e-21, 1.318912e-20, 5.080091e-21, -5.438722e-20, -5.920958e-21, 
    2.889679e-20, 3.004008e-21, -8.562225e-21, 3.154704e-21, 5.772229e-21, 
    -1.02326e-20, -3.080334e-21, -1.244835e-20, -2.153786e-20, 1.799887e-21, 
    -3.197486e-20, 2.410704e-20, 1.421203e-20, -1.879594e-20, -2.791259e-20, 
    -2.654263e-21, -2.220145e-20, -1.180983e-21, 2.272648e-20, -4.849686e-21, 
    1.740066e-20, 2.864937e-20, -2.829653e-20, -2.472084e-20, -2.641356e-20, 
    3.299665e-20, -1.15504e-20, 2.801436e-20, -2.338044e-20, 1.627794e-20, 
    -8.351316e-21, -3.031581e-20, -3.110377e-20, -3.640102e-20, 
    -2.061167e-22, 5.259499e-20, 1.617787e-20, -6.806458e-21, 2.537623e-20, 
    -2.1619e-20, -1.340852e-20, -3.391836e-20, 7.521782e-21, -9.969644e-21, 
    -1.153288e-20, -2.151071e-20, 7.313102e-21, 1.650101e-20, -3.881582e-20, 
    -8.33151e-21, 1.988163e-20, -4.902828e-21, -1.750007e-22, 2.282713e-20, 
    -3.386805e-20, 3.796962e-20, 1.366466e-20, -2.986005e-20, 8.277797e-21, 
    -3.072972e-20, -2.855294e-21, 6.027804e-21, -1.826129e-20, 4.48186e-21, 
    -3.833236e-20, 4.11868e-20, 3.064972e-20, -1.039572e-20, -2.478842e-20, 
    1.225326e-20, 8.213877e-21, 1.485497e-20, 1.954263e-20, -2.116241e-20, 
    3.879072e-21, -3.566988e-20, -1.709729e-20, -7.981783e-21, -2.017059e-20, 
    1.344356e-20, 2.647181e-20, -5.320936e-20, 2.832002e-20, -3.242214e-20, 
    -4.37031e-20, -2.13504e-20, 1.955819e-20, 1.74507e-20, -1.520866e-20, 
    3.408233e-20, 6.741687e-20, 8.750249e-21, 1.089022e-20, 1.938487e-20, 
    -3.552231e-21, -1.141467e-20, 2.29091e-20, 1.518717e-20, -1.231291e-21, 
    -7.011665e-22, -5.002913e-21, -1.759887e-20, 1.623553e-20, 5.878545e-21, 
    -5.419678e-21, -6.131295e-21, -3.788282e-20, 2.427442e-20, 3.120754e-20, 
    8.939096e-21, -1.543598e-20, 1.682956e-20, -7.673581e-21, -2.288902e-20, 
    7.861605e-21, 3.378885e-20, -6.756974e-21, -1.660563e-20, 2.564624e-20, 
    1.528783e-20, 1.246445e-20, -3.136756e-20, 7.258271e-21, -2.885266e-20, 
    -1.871253e-20, 3.159942e-20, 2.450993e-20, 7.297859e-21, 5.722331e-20, 
    1.495052e-20, -3.36659e-20, -4.268102e-20, -1.765033e-20, 1.607664e-20, 
    2.426366e-20, -1.594658e-20, 2.987419e-20, 1.831539e-21, -1.910684e-21, 
    4.010083e-20, -3.51587e-20, 1.173757e-20, -2.682437e-20, 4.92857e-21, 
    4.273306e-20, -1.374077e-21, -2.439994e-20, 3.391414e-20, -3.374109e-20, 
    1.122015e-20, -3.663879e-20, -6.293576e-21, 1.194679e-20, -2.603526e-20, 
    -1.301664e-20, -3.292541e-20, 2.431711e-20, -4.668717e-21, 2.248303e-20, 
    -2.948288e-20, -2.587413e-20, 8.466081e-21, 1.352867e-20, 1.324227e-20, 
    1.424679e-21, 6.714845e-21, -2.228764e-21, 1.917312e-20, 1.135134e-20, 
    7.283703e-21, 1.817675e-20, 6.477365e-21, 2.268064e-20, 6.12452e-21, 
    2.251389e-21, -2.966581e-20, -1.518207e-20, 1.257501e-20, 2.776389e-20, 
    2.54633e-20, 2.36476e-20, 3.339332e-20, -2.61051e-20, -2.740227e-20, 
    -1.229569e-20, -3.750983e-21, 1.513457e-20, 2.71399e-20, 1.67733e-20, 
    1.420498e-20, -3.026068e-20, 1.563416e-20, -2.45645e-20, -3.280541e-21, 
    -7.661145e-21, -8.530546e-21, 3.122592e-20, -3.534758e-20, -1.260889e-22, 
    -1.62067e-20, -1.809843e-20, 6.798269e-21, 2.576131e-20, -6.301503e-21, 
    -4.038525e-20, -3.690225e-21, -1.873287e-20, -2.005041e-20, 9.01798e-21, 
    -1.082321e-20, 2.276917e-20, -3.246825e-20, -2.282285e-20, 1.933597e-20, 
    -4.545452e-21, -1.992912e-20, -1.896587e-20, -3.356002e-21, 8.5755e-21, 
    -4.195075e-20, 1.303898e-20, 4.981603e-20, 1.796416e-20, 2.269877e-20, 
    -2.191501e-20, 3.894887e-21, -8.708692e-21, -2.541552e-20, 8.931186e-21, 
    -3.441627e-20, 8.381833e-21, -1.008303e-20, 1.794575e-20, -1.157783e-20, 
    8.412647e-21, 2.429337e-20, -2.107985e-20, -8.766347e-21, 3.375834e-20, 
    -3.246314e-20, 1.488097e-20, -2.158677e-20, -7.465522e-21, -1.496325e-20, 
    8.387787e-21, 4.224131e-22, 9.440393e-21, -1.392455e-21, 1.086676e-20, 
    -1.025041e-20, 1.871141e-20, 5.593544e-21, -1.491799e-20, 5.220926e-21 ;

 M_SOIL2C_TO_LEACHING =
  3.643155e-20, 4.356713e-20, 8.282883e-21, 8.587657e-21, 7.398778e-21, 
    2.282599e-20, -1.348343e-20, 1.379838e-20, -2.652863e-20, 2.503017e-20, 
    3.614133e-21, -2.518396e-20, 1.665844e-21, -2.423004e-20, 1.087977e-20, 
    -4.938825e-20, -1.186736e-20, 2.042448e-21, -1.532599e-20, -1.761979e-20, 
    -1.576762e-20, 3.547027e-20, 2.620333e-21, 2.841741e-21, -2.319233e-21, 
    5.056644e-21, 1.714224e-20, 2.23346e-20, -1.766248e-20, -5.99558e-21, 
    8.268725e-21, -6.182468e-21, -2.03651e-20, 1.9904e-20, -9.463e-21, 
    3.73674e-20, 3.21858e-21, 6.238625e-20, 6.00181e-21, -1.897774e-20, 
    2.0144e-20, 2.68617e-20, -5.918124e-21, 2.295519e-20, 1.998229e-20, 
    7.693413e-21, 1.710797e-21, 3.359547e-20, 3.05065e-21, 1.101491e-20, 
    3.465684e-20, -2.567958e-20, 2.123619e-20, -1.089649e-21, 5.39085e-21, 
    1.359933e-20, 6.746524e-21, 4.037932e-20, -6.206799e-21, 1.375795e-20, 
    -4.592932e-20, -3.520268e-21, 1.130062e-21, 5.010278e-21, -1.151273e-21, 
    1.545436e-20, 1.272542e-20, 1.871789e-20, 9.396845e-21, 1.948073e-20, 
    -1.321852e-20, 1.880979e-20, 1.34707e-20, -2.044626e-20, -2.922673e-20, 
    -8.061212e-21, 2.926885e-20, 2.57853e-22, -7.178252e-21, -1.324395e-20, 
    -1.538818e-20, -4.269461e-20, -1.000189e-20, -3.439957e-20, -1.03259e-20, 
    -2.063031e-20, -2.910007e-20, -2.47135e-20, -3.782933e-22, -1.724232e-20, 
    1.527282e-20, -2.637144e-20, -2.513844e-20, -4.085492e-22, 2.646163e-20, 
    2.42549e-20, -1.886181e-20, -8.480801e-21, 3.852785e-21, 1.004287e-20, 
    -9.833333e-22, -1.615327e-20, -1.108598e-21, 5.457839e-21, -6.775923e-21, 
    -3.272032e-21, -3.769933e-21, 1.862122e-20, 1.011836e-20, 4.208454e-21, 
    -5.074181e-21, 1.080088e-20, 3.87651e-21, 7.100765e-21, -1.66749e-20, 
    -1.065754e-20, -2.118501e-20, -1.143562e-20, -2.035949e-21, -3.49187e-22, 
    3.146936e-20, 2.164444e-20, -1.48951e-20, -1.073642e-20, -6.794017e-21, 
    -1.11147e-20, -2.94645e-20, 8.121452e-21, 1.249247e-20, -5.713134e-21, 
    -8.315123e-21, 1.999556e-20, -4.86721e-20, -2.43598e-20, 1.50509e-20, 
    2.685208e-20, 3.255934e-21, -2.996374e-21, -6.515809e-21, 2.421052e-20, 
    -2.445396e-20, -2.294586e-20, -1.066093e-20, -3.151046e-21, 1.322218e-20, 
    1.097419e-20, 2.463828e-20, 2.100861e-20, 2.600982e-20, -2.850887e-20, 
    3.784238e-20, -4.53612e-21, -2.901927e-21, -6.91356e-20, -5.248701e-20, 
    -7.855956e-21, 4.712863e-21, -1.682515e-21, -4.945726e-20, 2.5149e-21, 
    -2.662452e-21, -3.626925e-20, -1.140139e-20, -2.895049e-20, 
    -5.153343e-21, -1.345912e-20, 1.083083e-20, -1.673315e-20, -2.426423e-20, 
    -2.375816e-20, -8.60362e-22, -3.183353e-20, 1.385605e-20, -6.063734e-21, 
    -2.342847e-20, -1.269122e-20, 1.001376e-20, 4.897464e-21, 2.380509e-20, 
    -6.170622e-21, -2.450174e-20, 5.389117e-21, -2.690579e-20, -8.987178e-21, 
    -5.585289e-20, 3.978874e-21, -9.677306e-21, -2.428516e-20, 1.168976e-20, 
    7.379274e-21, 5.220311e-20, 2.65719e-20, 1.283287e-20, -1.151872e-20, 
    1.222555e-20, 1.505543e-20, -1.426857e-20, -2.639347e-20, 1.195864e-20, 
    -1.436894e-20, 2.197017e-20, 6.042533e-21, -6.762649e-21, -3.196866e-20, 
    7.17314e-21, -4.509553e-21, 1.240906e-20, 2.864089e-20, -1.729067e-20, 
    3.718617e-20, -4.988079e-20, 1.014239e-20, 2.411326e-20, 3.147445e-20, 
    4.971058e-20, -3.133023e-20, -2.061504e-20, 5.087455e-21, 2.446809e-20, 
    1.300958e-20, 2.75049e-20, -1.429796e-20, -1.476307e-20, 2.443659e-21, 
    -9.610579e-21, -2.536917e-20, -1.54371e-20, 4.634498e-21, 9.81952e-21, 
    2.128228e-20, 8.277797e-21, 6.311954e-21, -1.497888e-21, 2.564735e-20, 
    1.248115e-20, 4.079793e-21, -9.344215e-22, -1.128777e-20, -1.792431e-20, 
    2.566291e-20, -1.414079e-20, 1.106891e-20, -1.837384e-20, 8.444046e-21, 
    -1.089473e-20, 4.338511e-21, 5.706044e-20, 3.904371e-20, -4.43794e-20, 
    3.178431e-20, 2.18285e-20, -2.42473e-20, -1.730114e-20, -4.280684e-20, 
    8.640537e-21, 3.238735e-20, 3.22058e-21, 2.650322e-21, 7.111526e-21, 
    5.216957e-21, 4.124484e-21, 2.836345e-21, -1.900885e-20, -1.960907e-20, 
    -3.506541e-20, -1.253637e-21, 6.795445e-21, 3.041787e-20, -2.845147e-20, 
    4.960059e-20, -2.819958e-21, 1.400959e-20, 1.563556e-20, -1.484901e-20, 
    1.837298e-20, -1.281788e-20, -1.108783e-20, 4.031996e-20, 1.417641e-20, 
    1.174379e-20, -1.16618e-20, -2.346943e-21, -2.243865e-20, -6.067964e-21, 
    -1.127503e-20, 6.448804e-21, -1.378735e-20, 2.41664e-20, 4.911883e-20, 
    -1.897154e-20, 3.73712e-21, -1.149583e-21, 1.262901e-20, 1.514927e-20, 
    3.090304e-20, 5.198543e-20, 1.771902e-20, -3.197261e-20, 6.42083e-22, 
    -3.809825e-20, -3.994929e-20, 2.083953e-20, 3.23416e-21, 2.516049e-20, 
    -2.518396e-20, 1.001434e-20, -3.079216e-21, -7.15932e-21, -5.377965e-20, 
    4.442255e-21, 1.57054e-20, -8.831384e-21, 1.056846e-20, -5.336065e-20, 
    4.083649e-20, 2.022034e-20, -2.47788e-20, -2.906489e-22, -3.087591e-20, 
    2.166736e-20, -2.417659e-20, -1.932154e-20, -7.316498e-21, 5.604567e-21, 
    7.878302e-21, 1.502036e-20, 2.502336e-20, -7.832776e-21, -4.492705e-20, 
    5.211831e-20, 3.494354e-20, -6.060051e-20, 5.522524e-20, 5.076515e-20, 
    1.444811e-20, -2.199135e-20, -1.609813e-20, 2.041655e-20 ;

 M_SOIL3C_TO_LEACHING =
  1.374834e-20, 4.872578e-21, -2.790977e-20, -1.127982e-20, -2.075612e-20, 
    -1.875919e-20, -4.464659e-20, 2.456362e-21, 2.280082e-20, -2.089637e-20, 
    3.03028e-20, -1.886407e-20, -1.511477e-20, 2.379168e-21, -5.184995e-21, 
    1.807513e-21, 2.393031e-21, 2.567564e-20, 2.117765e-20, -7.9142e-21, 
    9.944213e-21, -3.14965e-20, -3.236133e-21, 1.509783e-21, -1.699945e-20, 
    -4.101433e-20, 1.059115e-21, -1.528697e-20, -2.391704e-20, 2.970933e-21, 
    -4.948377e-23, -1.774954e-20, -2.962623e-20, -4.717629e-21, 
    -2.426226e-20, 2.459957e-20, -3.545515e-22, 1.356628e-20, 3.727833e-20, 
    5.301189e-21, -2.280527e-21, 9.808029e-22, -1.99721e-20, 3.248718e-20, 
    3.200428e-20, 9.914813e-21, -1.717335e-20, 3.315868e-21, 1.194282e-20, 
    3.002516e-20, -1.522196e-20, -1.602376e-20, -1.303475e-20, 2.862395e-20, 
    -1.282494e-20, 2.251357e-20, -2.265211e-20, 1.456629e-20, 1.451849e-20, 
    1.822494e-21, 9.236253e-21, 9.232858e-21, -2.396822e-20, 1.703904e-20, 
    -1.847533e-20, -7.230822e-21, 3.675134e-20, 3.96431e-20, -1.8872e-20, 
    4.491658e-20, 3.171532e-20, -1.021506e-20, 1.83481e-20, -2.839099e-20, 
    3.152081e-20, 1.41074e-20, -2.087288e-20, -3.877598e-20, 3.315296e-21, 
    -2.676037e-21, -9.77317e-21, 1.916265e-20, -1.69073e-21, -3.768798e-21, 
    1.062728e-20, -3.228106e-20, -4.732903e-21, 1.91408e-21, 6.467181e-21, 
    -6.949244e-21, 2.23776e-20, -7.272117e-21, 5.639632e-21, 3.017593e-21, 
    8.105898e-21, 2.103526e-21, 1.29273e-20, 2.07072e-20, -2.935679e-20, 
    -1.347693e-20, -3.13195e-20, 2.229043e-21, 1.070702e-20, 1.830737e-20, 
    2.234027e-20, -4.699251e-21, 2.612205e-20, 1.015795e-20, 2.195113e-21, 
    2.181069e-20, 2.677405e-20, 3.269386e-20, -2.051635e-20, -4.231971e-20, 
    7.400175e-21, 3.636371e-20, 1.822144e-20, -1.229229e-20, -1.252101e-20, 
    -1.156935e-20, -6.132723e-21, 8.397387e-21, -1.322273e-20, 8.91053e-21, 
    -2.455346e-20, 1.394145e-21, -1.22117e-20, 2.438044e-20, 1.692002e-20, 
    2.763666e-20, -4.279973e-21, 3.320399e-21, -1.638412e-21, -8.162441e-21, 
    -2.647096e-20, -2.396765e-20, 5.657447e-21, 3.407473e-20, 5.374987e-21, 
    -5.419939e-21, 2.083726e-21, 6.719386e-21, 2.272251e-20, -5.317064e-20, 
    -1.946432e-20, -3.884437e-21, 1.177856e-21, 2.191587e-20, -3.432465e-20, 
    -4.219467e-21, 4.916103e-21, -3.348775e-20, 4.54863e-20, 2.179685e-20, 
    4.071214e-22, -1.36573e-20, 4.729916e-20, 1.004599e-20, 1.643938e-20, 
    2.126729e-20, -1.538932e-20, 3.157707e-20, -5.51291e-20, -2.966496e-20, 
    3.519445e-21, -1.139715e-20, -6.972136e-21, -7.991116e-21, -2.465782e-20, 
    2.044512e-20, -1.715217e-20, -4.950107e-20, -3.414682e-20, -2.903195e-20, 
    4.199399e-20, 2.742207e-20, -3.799905e-21, -1.520752e-20, 1.247946e-20, 
    -2.05155e-20, -3.150736e-21, 1.270225e-20, 8.815269e-21, -2.003486e-20, 
    -8.890201e-21, -6.931723e-21, -3.713443e-20, 3.551805e-20, 1.757341e-20, 
    2.021443e-20, 9.615664e-21, 4.430522e-22, -3.996146e-20, -1.245572e-20, 
    -1.693558e-20, 3.136191e-20, -1.098212e-20, -1.668224e-20, -5.52535e-20, 
    -9.648478e-21, -3.146003e-20, 4.526375e-23, 1.108812e-20, 1.508822e-20, 
    4.094496e-21, -1.491999e-20, 1.148e-20, 1.823189e-20, -4.232741e-21, 
    2.18073e-20, 1.007398e-20, -4.350096e-21, 3.080861e-20, -3.560315e-20, 
    2.175755e-20, -2.822473e-20, 2.287582e-21, 1.290071e-20, -4.396557e-22, 
    9.950711e-21, 2.071425e-20, 2.524886e-22, -2.425038e-20, 2.633079e-21, 
    2.098795e-20, 3.68811e-20, -1.874249e-20, -4.641569e-21, -2.137104e-20, 
    1.939194e-20, -7.174023e-21, 1.427139e-20, 5.172838e-21, 4.031737e-21, 
    -1.83362e-20, 1.342067e-20, -2.254636e-20, -1.552985e-20, 2.450653e-20, 
    2.726796e-20, 2.133345e-20, -3.110831e-20, -2.145842e-20, -2.52535e-21, 
    -1.709786e-20, 4.402977e-21, 3.115409e-21, -5.230322e-20, 3.997513e-21, 
    4.127164e-20, -1.176555e-20, 1.001122e-20, -1.838881e-20, -6.060338e-21, 
    -1.563868e-20, -1.871084e-20, 1.826245e-20, 2.114539e-21, 3.02047e-20, 
    9.823462e-21, 2.018641e-20, 7.394004e-21, 2.220736e-20, 1.852847e-20, 
    -1.189959e-20, -1.920873e-21, -5.766408e-20, -7.930325e-21, 
    -1.400448e-20, -2.345307e-20, 1.152043e-20, 1.54162e-20, -2.005609e-20, 
    -1.427649e-20, 2.445396e-20, -3.907764e-20, -2.751933e-20, -1.721858e-20, 
    5.405671e-20, 3.033305e-20, 2.533605e-20, -8.942208e-21, 3.650898e-21, 
    -1.094873e-20, -3.409111e-20, 5.483009e-21, 2.599991e-20, 2.040328e-20, 
    -1.48677e-20, -1.236607e-20, 1.387303e-20, 2.456167e-20, -1.096374e-20, 
    1.039685e-20, 2.219407e-20, -6.639384e-21, 1.479249e-21, -9.15568e-21, 
    4.471811e-20, 3.969088e-20, 1.605966e-20, -6.741421e-21, 2.028818e-20, 
    1.156822e-20, 1.820785e-20, -1.151845e-21, 5.162388e-21, -1.473196e-20, 
    -1.733111e-20, -1.71445e-20, 2.807093e-20, 1.403108e-20, -1.34464e-20, 
    -3.913265e-21, -6.803061e-21, 4.831981e-20, 1.272345e-20, 2.637593e-21, 
    5.222616e-21, -1.002336e-20, -1.245542e-20, 1.653687e-21, 1.131516e-21, 
    -7.324998e-21, 3.395036e-21, -4.055479e-21, -4.623015e-20, 1.709898e-20, 
    -1.798959e-20, -1.868427e-20, -5.286217e-20, 3.282392e-20, 3.290928e-20, 
    1.156935e-20, -2.405278e-20, 3.941521e-20, 2.011489e-20, 2.469683e-20 ;

 NBP =
  -7.623649e-08, -7.644516e-08, -7.640461e-08, -7.657286e-08, -7.647954e-08, 
    -7.658971e-08, -7.627882e-08, -7.645342e-08, -7.634197e-08, -7.62553e-08, 
    -7.689925e-08, -7.658038e-08, -7.723048e-08, -7.70272e-08, -7.753781e-08, 
    -7.719884e-08, -7.760615e-08, -7.752807e-08, -7.776314e-08, -7.76958e-08, 
    -7.799632e-08, -7.779421e-08, -7.815211e-08, -7.794808e-08, 
    -7.797998e-08, -7.778754e-08, -7.664459e-08, -7.685954e-08, 
    -7.663184e-08, -7.66625e-08, -7.664875e-08, -7.648146e-08, -7.639712e-08, 
    -7.622056e-08, -7.625263e-08, -7.638231e-08, -7.667629e-08, 
    -7.657653e-08, -7.682798e-08, -7.682231e-08, -7.710213e-08, 
    -7.697598e-08, -7.744618e-08, -7.731258e-08, -7.769862e-08, 
    -7.760154e-08, -7.769405e-08, -7.766601e-08, -7.769442e-08, 
    -7.755205e-08, -7.761304e-08, -7.748777e-08, -7.69996e-08, -7.714308e-08, 
    -7.671504e-08, -7.64575e-08, -7.628647e-08, -7.616506e-08, -7.618222e-08, 
    -7.621494e-08, -7.638307e-08, -7.654115e-08, -7.666159e-08, 
    -7.674213e-08, -7.682149e-08, -7.706157e-08, -7.718869e-08, 
    -7.747317e-08, -7.742187e-08, -7.750881e-08, -7.759189e-08, 
    -7.773131e-08, -7.770838e-08, -7.776979e-08, -7.750653e-08, 
    -7.768149e-08, -7.739264e-08, -7.747165e-08, -7.684295e-08, 
    -7.660345e-08, -7.650154e-08, -7.64124e-08, -7.619542e-08, -7.634526e-08, 
    -7.628619e-08, -7.642673e-08, -7.651601e-08, -7.647186e-08, 
    -7.674434e-08, -7.663841e-08, -7.719622e-08, -7.695601e-08, 
    -7.758219e-08, -7.74324e-08, -7.76181e-08, -7.752336e-08, -7.768568e-08, 
    -7.75396e-08, -7.779266e-08, -7.784774e-08, -7.781009e-08, -7.795472e-08, 
    -7.753149e-08, -7.769404e-08, -7.647062e-08, -7.647782e-08, 
    -7.651137e-08, -7.636387e-08, -7.635484e-08, -7.621968e-08, 
    -7.633997e-08, -7.639117e-08, -7.65212e-08, -7.659807e-08, -7.667116e-08, 
    -7.683181e-08, -7.701119e-08, -7.726197e-08, -7.744212e-08, 
    -7.756284e-08, -7.748882e-08, -7.755416e-08, -7.748111e-08, 
    -7.744688e-08, -7.782709e-08, -7.761361e-08, -7.793392e-08, 
    -7.791621e-08, -7.777125e-08, -7.791819e-08, -7.648288e-08, 
    -7.644144e-08, -7.629752e-08, -7.641015e-08, -7.620496e-08, 
    -7.631981e-08, -7.638584e-08, -7.66406e-08, -7.669659e-08, -7.674847e-08, 
    -7.685095e-08, -7.698243e-08, -7.721304e-08, -7.741363e-08, 
    -7.759672e-08, -7.758331e-08, -7.758803e-08, -7.762892e-08, 
    -7.752763e-08, -7.764555e-08, -7.766533e-08, -7.76136e-08, -7.791383e-08, 
    -7.782807e-08, -7.791583e-08, -7.785999e-08, -7.645492e-08, 
    -7.652464e-08, -7.648696e-08, -7.65578e-08, -7.650789e-08, -7.672979e-08, 
    -7.679631e-08, -7.710752e-08, -7.697984e-08, -7.718307e-08, 
    -7.700049e-08, -7.703284e-08, -7.718965e-08, -7.701037e-08, 
    -7.740255e-08, -7.713665e-08, -7.76305e-08, -7.736501e-08, -7.764714e-08, 
    -7.759594e-08, -7.768072e-08, -7.775665e-08, -7.785217e-08, 
    -7.802836e-08, -7.798757e-08, -7.813491e-08, -7.662858e-08, 
    -7.671898e-08, -7.671105e-08, -7.680566e-08, -7.687562e-08, 
    -7.702726e-08, -7.727039e-08, -7.717897e-08, -7.73468e-08, -7.738048e-08, 
    -7.712552e-08, -7.728205e-08, -7.67795e-08, -7.686069e-08, -7.681236e-08, 
    -7.66357e-08, -7.720001e-08, -7.691045e-08, -7.744509e-08, -7.728828e-08, 
    -7.774582e-08, -7.751829e-08, -7.796511e-08, -7.815598e-08, 
    -7.833569e-08, -7.854553e-08, -7.676834e-08, -7.670692e-08, 
    -7.681692e-08, -7.696904e-08, -7.711023e-08, -7.729785e-08, 
    -7.731705e-08, -7.735219e-08, -7.744323e-08, -7.751974e-08, 
    -7.736328e-08, -7.753892e-08, -7.687949e-08, -7.722515e-08, 
    -7.668368e-08, -7.684673e-08, -7.696008e-08, -7.691038e-08, 
    -7.716854e-08, -7.722935e-08, -7.747646e-08, -7.734874e-08, 
    -7.810886e-08, -7.777265e-08, -7.870533e-08, -7.844478e-08, 
    -7.668545e-08, -7.676814e-08, -7.705584e-08, -7.691897e-08, 
    -7.731038e-08, -7.740669e-08, -7.748498e-08, -7.758503e-08, 
    -7.759585e-08, -7.765512e-08, -7.755798e-08, -7.765129e-08, 
    -7.729825e-08, -7.745604e-08, -7.702298e-08, -7.71284e-08, -7.707991e-08, 
    -7.702671e-08, -7.71909e-08, -7.736573e-08, -7.736951e-08, -7.742555e-08, 
    -7.758342e-08, -7.731197e-08, -7.815218e-08, -7.763335e-08, -7.68583e-08, 
    -7.701748e-08, -7.704026e-08, -7.697859e-08, -7.739703e-08, 
    -7.724544e-08, -7.765367e-08, -7.754338e-08, -7.77241e-08, -7.76343e-08, 
    -7.762108e-08, -7.750573e-08, -7.74339e-08, -7.725239e-08, -7.710467e-08, 
    -7.698755e-08, -7.701478e-08, -7.714345e-08, -7.737644e-08, 
    -7.759681e-08, -7.754854e-08, -7.771037e-08, -7.728201e-08, 
    -7.746164e-08, -7.739221e-08, -7.757325e-08, -7.717654e-08, 
    -7.751427e-08, -7.709018e-08, -7.712737e-08, -7.724243e-08, -7.74738e-08, 
    -7.752503e-08, -7.757966e-08, -7.754596e-08, -7.738236e-08, 
    -7.735557e-08, -7.723964e-08, -7.720762e-08, -7.711928e-08, 
    -7.704612e-08, -7.711296e-08, -7.718313e-08, -7.738244e-08, -7.7562e-08, 
    -7.775772e-08, -7.780563e-08, -7.803415e-08, -7.784809e-08, 
    -7.815506e-08, -7.789401e-08, -7.834588e-08, -7.753389e-08, 
    -7.788639e-08, -7.724768e-08, -7.731652e-08, -7.744099e-08, 
    -7.772646e-08, -7.757239e-08, -7.775259e-08, -7.735452e-08, 
    -7.714787e-08, -7.709443e-08, -7.699466e-08, -7.709671e-08, 
    -7.708842e-08, -7.718606e-08, -7.715469e-08, -7.738906e-08, 
    -7.726317e-08, -7.762075e-08, -7.775118e-08, -7.811946e-08, 
    -7.834512e-08, -7.857481e-08, -7.867618e-08, -7.870703e-08, -7.871993e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  7.623649e-08, 7.644516e-08, 7.640461e-08, 7.657286e-08, 7.647954e-08, 
    7.658971e-08, 7.627882e-08, 7.645342e-08, 7.634197e-08, 7.62553e-08, 
    7.689925e-08, 7.658038e-08, 7.723048e-08, 7.70272e-08, 7.753781e-08, 
    7.719884e-08, 7.760615e-08, 7.752807e-08, 7.776314e-08, 7.76958e-08, 
    7.799632e-08, 7.779421e-08, 7.815211e-08, 7.794808e-08, 7.797998e-08, 
    7.778754e-08, 7.664459e-08, 7.685954e-08, 7.663184e-08, 7.66625e-08, 
    7.664875e-08, 7.648146e-08, 7.639712e-08, 7.622056e-08, 7.625263e-08, 
    7.638231e-08, 7.667629e-08, 7.657653e-08, 7.682798e-08, 7.682231e-08, 
    7.710213e-08, 7.697598e-08, 7.744618e-08, 7.731258e-08, 7.769862e-08, 
    7.760154e-08, 7.769405e-08, 7.766601e-08, 7.769442e-08, 7.755205e-08, 
    7.761304e-08, 7.748777e-08, 7.69996e-08, 7.714308e-08, 7.671504e-08, 
    7.64575e-08, 7.628647e-08, 7.616506e-08, 7.618222e-08, 7.621494e-08, 
    7.638307e-08, 7.654115e-08, 7.666159e-08, 7.674213e-08, 7.682149e-08, 
    7.706157e-08, 7.718869e-08, 7.747317e-08, 7.742187e-08, 7.750881e-08, 
    7.759189e-08, 7.773131e-08, 7.770838e-08, 7.776979e-08, 7.750653e-08, 
    7.768149e-08, 7.739264e-08, 7.747165e-08, 7.684295e-08, 7.660345e-08, 
    7.650154e-08, 7.64124e-08, 7.619542e-08, 7.634526e-08, 7.628619e-08, 
    7.642673e-08, 7.651601e-08, 7.647186e-08, 7.674434e-08, 7.663841e-08, 
    7.719622e-08, 7.695601e-08, 7.758219e-08, 7.74324e-08, 7.76181e-08, 
    7.752336e-08, 7.768568e-08, 7.75396e-08, 7.779266e-08, 7.784774e-08, 
    7.781009e-08, 7.795472e-08, 7.753149e-08, 7.769404e-08, 7.647062e-08, 
    7.647782e-08, 7.651137e-08, 7.636387e-08, 7.635484e-08, 7.621968e-08, 
    7.633997e-08, 7.639117e-08, 7.65212e-08, 7.659807e-08, 7.667116e-08, 
    7.683181e-08, 7.701119e-08, 7.726197e-08, 7.744212e-08, 7.756284e-08, 
    7.748882e-08, 7.755416e-08, 7.748111e-08, 7.744688e-08, 7.782709e-08, 
    7.761361e-08, 7.793392e-08, 7.791621e-08, 7.777125e-08, 7.791819e-08, 
    7.648288e-08, 7.644144e-08, 7.629752e-08, 7.641015e-08, 7.620496e-08, 
    7.631981e-08, 7.638584e-08, 7.66406e-08, 7.669659e-08, 7.674847e-08, 
    7.685095e-08, 7.698243e-08, 7.721304e-08, 7.741363e-08, 7.759672e-08, 
    7.758331e-08, 7.758803e-08, 7.762892e-08, 7.752763e-08, 7.764555e-08, 
    7.766533e-08, 7.76136e-08, 7.791383e-08, 7.782807e-08, 7.791583e-08, 
    7.785999e-08, 7.645492e-08, 7.652464e-08, 7.648696e-08, 7.65578e-08, 
    7.650789e-08, 7.672979e-08, 7.679631e-08, 7.710752e-08, 7.697984e-08, 
    7.718307e-08, 7.700049e-08, 7.703284e-08, 7.718965e-08, 7.701037e-08, 
    7.740255e-08, 7.713665e-08, 7.76305e-08, 7.736501e-08, 7.764714e-08, 
    7.759594e-08, 7.768072e-08, 7.775665e-08, 7.785217e-08, 7.802836e-08, 
    7.798757e-08, 7.813491e-08, 7.662858e-08, 7.671898e-08, 7.671105e-08, 
    7.680566e-08, 7.687562e-08, 7.702726e-08, 7.727039e-08, 7.717897e-08, 
    7.73468e-08, 7.738048e-08, 7.712552e-08, 7.728205e-08, 7.67795e-08, 
    7.686069e-08, 7.681236e-08, 7.66357e-08, 7.720001e-08, 7.691045e-08, 
    7.744509e-08, 7.728828e-08, 7.774582e-08, 7.751829e-08, 7.796511e-08, 
    7.815598e-08, 7.833569e-08, 7.854553e-08, 7.676834e-08, 7.670692e-08, 
    7.681692e-08, 7.696904e-08, 7.711023e-08, 7.729785e-08, 7.731705e-08, 
    7.735219e-08, 7.744323e-08, 7.751974e-08, 7.736328e-08, 7.753892e-08, 
    7.687949e-08, 7.722515e-08, 7.668368e-08, 7.684673e-08, 7.696008e-08, 
    7.691038e-08, 7.716854e-08, 7.722935e-08, 7.747646e-08, 7.734874e-08, 
    7.810886e-08, 7.777265e-08, 7.870533e-08, 7.844478e-08, 7.668545e-08, 
    7.676814e-08, 7.705584e-08, 7.691897e-08, 7.731038e-08, 7.740669e-08, 
    7.748498e-08, 7.758503e-08, 7.759585e-08, 7.765512e-08, 7.755798e-08, 
    7.765129e-08, 7.729825e-08, 7.745604e-08, 7.702298e-08, 7.71284e-08, 
    7.707991e-08, 7.702671e-08, 7.71909e-08, 7.736573e-08, 7.736951e-08, 
    7.742555e-08, 7.758342e-08, 7.731197e-08, 7.815218e-08, 7.763335e-08, 
    7.68583e-08, 7.701748e-08, 7.704026e-08, 7.697859e-08, 7.739703e-08, 
    7.724544e-08, 7.765367e-08, 7.754338e-08, 7.77241e-08, 7.76343e-08, 
    7.762108e-08, 7.750573e-08, 7.74339e-08, 7.725239e-08, 7.710467e-08, 
    7.698755e-08, 7.701478e-08, 7.714345e-08, 7.737644e-08, 7.759681e-08, 
    7.754854e-08, 7.771037e-08, 7.728201e-08, 7.746164e-08, 7.739221e-08, 
    7.757325e-08, 7.717654e-08, 7.751427e-08, 7.709018e-08, 7.712737e-08, 
    7.724243e-08, 7.74738e-08, 7.752503e-08, 7.757966e-08, 7.754596e-08, 
    7.738236e-08, 7.735557e-08, 7.723964e-08, 7.720762e-08, 7.711928e-08, 
    7.704612e-08, 7.711296e-08, 7.718313e-08, 7.738244e-08, 7.7562e-08, 
    7.775772e-08, 7.780563e-08, 7.803415e-08, 7.784809e-08, 7.815506e-08, 
    7.789401e-08, 7.834588e-08, 7.753389e-08, 7.788639e-08, 7.724768e-08, 
    7.731652e-08, 7.744099e-08, 7.772646e-08, 7.757239e-08, 7.775259e-08, 
    7.735452e-08, 7.714787e-08, 7.709443e-08, 7.699466e-08, 7.709671e-08, 
    7.708842e-08, 7.718606e-08, 7.715469e-08, 7.738906e-08, 7.726317e-08, 
    7.762075e-08, 7.775118e-08, 7.811946e-08, 7.834512e-08, 7.857481e-08, 
    7.867618e-08, 7.870703e-08, 7.871993e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -7.623649e-08, -7.644516e-08, -7.640461e-08, -7.657286e-08, -7.647954e-08, 
    -7.658971e-08, -7.627882e-08, -7.645342e-08, -7.634197e-08, -7.62553e-08, 
    -7.689925e-08, -7.658038e-08, -7.723048e-08, -7.70272e-08, -7.753781e-08, 
    -7.719884e-08, -7.760615e-08, -7.752807e-08, -7.776314e-08, -7.76958e-08, 
    -7.799632e-08, -7.779421e-08, -7.815211e-08, -7.794808e-08, 
    -7.797998e-08, -7.778754e-08, -7.664459e-08, -7.685954e-08, 
    -7.663184e-08, -7.66625e-08, -7.664875e-08, -7.648146e-08, -7.639712e-08, 
    -7.622056e-08, -7.625263e-08, -7.638231e-08, -7.667629e-08, 
    -7.657653e-08, -7.682798e-08, -7.682231e-08, -7.710213e-08, 
    -7.697598e-08, -7.744618e-08, -7.731258e-08, -7.769862e-08, 
    -7.760154e-08, -7.769405e-08, -7.766601e-08, -7.769442e-08, 
    -7.755205e-08, -7.761304e-08, -7.748777e-08, -7.69996e-08, -7.714308e-08, 
    -7.671504e-08, -7.64575e-08, -7.628647e-08, -7.616506e-08, -7.618222e-08, 
    -7.621494e-08, -7.638307e-08, -7.654115e-08, -7.666159e-08, 
    -7.674213e-08, -7.682149e-08, -7.706157e-08, -7.718869e-08, 
    -7.747317e-08, -7.742187e-08, -7.750881e-08, -7.759189e-08, 
    -7.773131e-08, -7.770838e-08, -7.776979e-08, -7.750653e-08, 
    -7.768149e-08, -7.739264e-08, -7.747165e-08, -7.684295e-08, 
    -7.660345e-08, -7.650154e-08, -7.64124e-08, -7.619542e-08, -7.634526e-08, 
    -7.628619e-08, -7.642673e-08, -7.651601e-08, -7.647186e-08, 
    -7.674434e-08, -7.663841e-08, -7.719622e-08, -7.695601e-08, 
    -7.758219e-08, -7.74324e-08, -7.76181e-08, -7.752336e-08, -7.768568e-08, 
    -7.75396e-08, -7.779266e-08, -7.784774e-08, -7.781009e-08, -7.795472e-08, 
    -7.753149e-08, -7.769404e-08, -7.647062e-08, -7.647782e-08, 
    -7.651137e-08, -7.636387e-08, -7.635484e-08, -7.621968e-08, 
    -7.633997e-08, -7.639117e-08, -7.65212e-08, -7.659807e-08, -7.667116e-08, 
    -7.683181e-08, -7.701119e-08, -7.726197e-08, -7.744212e-08, 
    -7.756284e-08, -7.748882e-08, -7.755416e-08, -7.748111e-08, 
    -7.744688e-08, -7.782709e-08, -7.761361e-08, -7.793392e-08, 
    -7.791621e-08, -7.777125e-08, -7.791819e-08, -7.648288e-08, 
    -7.644144e-08, -7.629752e-08, -7.641015e-08, -7.620496e-08, 
    -7.631981e-08, -7.638584e-08, -7.66406e-08, -7.669659e-08, -7.674847e-08, 
    -7.685095e-08, -7.698243e-08, -7.721304e-08, -7.741363e-08, 
    -7.759672e-08, -7.758331e-08, -7.758803e-08, -7.762892e-08, 
    -7.752763e-08, -7.764555e-08, -7.766533e-08, -7.76136e-08, -7.791383e-08, 
    -7.782807e-08, -7.791583e-08, -7.785999e-08, -7.645492e-08, 
    -7.652464e-08, -7.648696e-08, -7.65578e-08, -7.650789e-08, -7.672979e-08, 
    -7.679631e-08, -7.710752e-08, -7.697984e-08, -7.718307e-08, 
    -7.700049e-08, -7.703284e-08, -7.718965e-08, -7.701037e-08, 
    -7.740255e-08, -7.713665e-08, -7.76305e-08, -7.736501e-08, -7.764714e-08, 
    -7.759594e-08, -7.768072e-08, -7.775665e-08, -7.785217e-08, 
    -7.802836e-08, -7.798757e-08, -7.813491e-08, -7.662858e-08, 
    -7.671898e-08, -7.671105e-08, -7.680566e-08, -7.687562e-08, 
    -7.702726e-08, -7.727039e-08, -7.717897e-08, -7.73468e-08, -7.738048e-08, 
    -7.712552e-08, -7.728205e-08, -7.67795e-08, -7.686069e-08, -7.681236e-08, 
    -7.66357e-08, -7.720001e-08, -7.691045e-08, -7.744509e-08, -7.728828e-08, 
    -7.774582e-08, -7.751829e-08, -7.796511e-08, -7.815598e-08, 
    -7.833569e-08, -7.854553e-08, -7.676834e-08, -7.670692e-08, 
    -7.681692e-08, -7.696904e-08, -7.711023e-08, -7.729785e-08, 
    -7.731705e-08, -7.735219e-08, -7.744323e-08, -7.751974e-08, 
    -7.736328e-08, -7.753892e-08, -7.687949e-08, -7.722515e-08, 
    -7.668368e-08, -7.684673e-08, -7.696008e-08, -7.691038e-08, 
    -7.716854e-08, -7.722935e-08, -7.747646e-08, -7.734874e-08, 
    -7.810886e-08, -7.777265e-08, -7.870533e-08, -7.844478e-08, 
    -7.668545e-08, -7.676814e-08, -7.705584e-08, -7.691897e-08, 
    -7.731038e-08, -7.740669e-08, -7.748498e-08, -7.758503e-08, 
    -7.759585e-08, -7.765512e-08, -7.755798e-08, -7.765129e-08, 
    -7.729825e-08, -7.745604e-08, -7.702298e-08, -7.71284e-08, -7.707991e-08, 
    -7.702671e-08, -7.71909e-08, -7.736573e-08, -7.736951e-08, -7.742555e-08, 
    -7.758342e-08, -7.731197e-08, -7.815218e-08, -7.763335e-08, -7.68583e-08, 
    -7.701748e-08, -7.704026e-08, -7.697859e-08, -7.739703e-08, 
    -7.724544e-08, -7.765367e-08, -7.754338e-08, -7.77241e-08, -7.76343e-08, 
    -7.762108e-08, -7.750573e-08, -7.74339e-08, -7.725239e-08, -7.710467e-08, 
    -7.698755e-08, -7.701478e-08, -7.714345e-08, -7.737644e-08, 
    -7.759681e-08, -7.754854e-08, -7.771037e-08, -7.728201e-08, 
    -7.746164e-08, -7.739221e-08, -7.757325e-08, -7.717654e-08, 
    -7.751427e-08, -7.709018e-08, -7.712737e-08, -7.724243e-08, -7.74738e-08, 
    -7.752503e-08, -7.757966e-08, -7.754596e-08, -7.738236e-08, 
    -7.735557e-08, -7.723964e-08, -7.720762e-08, -7.711928e-08, 
    -7.704612e-08, -7.711296e-08, -7.718313e-08, -7.738244e-08, -7.7562e-08, 
    -7.775772e-08, -7.780563e-08, -7.803415e-08, -7.784809e-08, 
    -7.815506e-08, -7.789401e-08, -7.834588e-08, -7.753389e-08, 
    -7.788639e-08, -7.724768e-08, -7.731652e-08, -7.744099e-08, 
    -7.772646e-08, -7.757239e-08, -7.775259e-08, -7.735452e-08, 
    -7.714787e-08, -7.709443e-08, -7.699466e-08, -7.709671e-08, 
    -7.708842e-08, -7.718606e-08, -7.715469e-08, -7.738906e-08, 
    -7.726317e-08, -7.762075e-08, -7.775118e-08, -7.811946e-08, 
    -7.834512e-08, -7.857481e-08, -7.867618e-08, -7.870703e-08, -7.871993e-08 ;

 NET_NMIN =
  1.074021e-08, 1.07696e-08, 1.076389e-08, 1.078759e-08, 1.077445e-08, 
    1.078996e-08, 1.074617e-08, 1.077077e-08, 1.075507e-08, 1.074286e-08, 
    1.083357e-08, 1.078865e-08, 1.088023e-08, 1.085159e-08, 1.092352e-08, 
    1.087577e-08, 1.093315e-08, 1.092215e-08, 1.095526e-08, 1.094577e-08, 
    1.098811e-08, 1.095964e-08, 1.101005e-08, 1.098131e-08, 1.098581e-08, 
    1.09587e-08, 1.079769e-08, 1.082797e-08, 1.07959e-08, 1.080022e-08, 
    1.079828e-08, 1.077472e-08, 1.076283e-08, 1.073796e-08, 1.074248e-08, 
    1.076075e-08, 1.080216e-08, 1.078811e-08, 1.082353e-08, 1.082273e-08, 
    1.086215e-08, 1.084438e-08, 1.091061e-08, 1.089179e-08, 1.094617e-08, 
    1.09325e-08, 1.094553e-08, 1.094158e-08, 1.094558e-08, 1.092552e-08, 
    1.093412e-08, 1.091647e-08, 1.08477e-08, 1.086792e-08, 1.080762e-08, 
    1.077134e-08, 1.074725e-08, 1.073014e-08, 1.073256e-08, 1.073717e-08, 
    1.076086e-08, 1.078312e-08, 1.080009e-08, 1.081143e-08, 1.082261e-08, 
    1.085643e-08, 1.087434e-08, 1.091441e-08, 1.090719e-08, 1.091943e-08, 
    1.093114e-08, 1.095078e-08, 1.094755e-08, 1.09562e-08, 1.091911e-08, 
    1.094376e-08, 1.090307e-08, 1.09142e-08, 1.082564e-08, 1.07919e-08, 
    1.077754e-08, 1.076499e-08, 1.073442e-08, 1.075553e-08, 1.074721e-08, 
    1.076701e-08, 1.077958e-08, 1.077336e-08, 1.081174e-08, 1.079682e-08, 
    1.08754e-08, 1.084156e-08, 1.092977e-08, 1.090867e-08, 1.093483e-08, 
    1.092148e-08, 1.094435e-08, 1.092377e-08, 1.095942e-08, 1.096718e-08, 
    1.096187e-08, 1.098225e-08, 1.092263e-08, 1.094553e-08, 1.077319e-08, 
    1.07742e-08, 1.077893e-08, 1.075815e-08, 1.075688e-08, 1.073784e-08, 
    1.075478e-08, 1.0762e-08, 1.078031e-08, 1.079114e-08, 1.080144e-08, 
    1.082407e-08, 1.084934e-08, 1.088466e-08, 1.091004e-08, 1.092704e-08, 
    1.091662e-08, 1.092582e-08, 1.091553e-08, 1.091071e-08, 1.096427e-08, 
    1.09342e-08, 1.097932e-08, 1.097682e-08, 1.09564e-08, 1.09771e-08, 
    1.077491e-08, 1.076908e-08, 1.07488e-08, 1.076467e-08, 1.073576e-08, 
    1.075194e-08, 1.076124e-08, 1.079713e-08, 1.080502e-08, 1.081233e-08, 
    1.082676e-08, 1.084528e-08, 1.087777e-08, 1.090603e-08, 1.093182e-08, 
    1.092993e-08, 1.093059e-08, 1.093635e-08, 1.092208e-08, 1.09387e-08, 
    1.094148e-08, 1.093419e-08, 1.097649e-08, 1.096441e-08, 1.097677e-08, 
    1.09689e-08, 1.077098e-08, 1.07808e-08, 1.077549e-08, 1.078547e-08, 
    1.077844e-08, 1.08097e-08, 1.081907e-08, 1.086291e-08, 1.084492e-08, 
    1.087355e-08, 1.084783e-08, 1.085239e-08, 1.087447e-08, 1.084922e-08, 
    1.090446e-08, 1.086701e-08, 1.093658e-08, 1.089918e-08, 1.093892e-08, 
    1.093171e-08, 1.094365e-08, 1.095434e-08, 1.09678e-08, 1.099262e-08, 
    1.098687e-08, 1.100763e-08, 1.079544e-08, 1.080817e-08, 1.080706e-08, 
    1.082038e-08, 1.083024e-08, 1.08516e-08, 1.088585e-08, 1.087297e-08, 
    1.089661e-08, 1.090136e-08, 1.086544e-08, 1.088749e-08, 1.08167e-08, 
    1.082814e-08, 1.082133e-08, 1.079644e-08, 1.087593e-08, 1.083514e-08, 
    1.091046e-08, 1.088837e-08, 1.095282e-08, 1.092077e-08, 1.098371e-08, 
    1.10106e-08, 1.103591e-08, 1.106547e-08, 1.081513e-08, 1.080647e-08, 
    1.082197e-08, 1.08434e-08, 1.086329e-08, 1.088972e-08, 1.089242e-08, 
    1.089737e-08, 1.091019e-08, 1.092097e-08, 1.089893e-08, 1.092368e-08, 
    1.083078e-08, 1.087948e-08, 1.08032e-08, 1.082617e-08, 1.084214e-08, 
    1.083514e-08, 1.08715e-08, 1.088007e-08, 1.091488e-08, 1.089689e-08, 
    1.100396e-08, 1.09566e-08, 1.108798e-08, 1.105128e-08, 1.080345e-08, 
    1.08151e-08, 1.085562e-08, 1.083635e-08, 1.089148e-08, 1.090505e-08, 
    1.091608e-08, 1.093017e-08, 1.093169e-08, 1.094004e-08, 1.092636e-08, 
    1.09395e-08, 1.088977e-08, 1.0912e-08, 1.0851e-08, 1.086585e-08, 
    1.085902e-08, 1.085152e-08, 1.087465e-08, 1.089928e-08, 1.089981e-08, 
    1.090771e-08, 1.092994e-08, 1.089171e-08, 1.101006e-08, 1.093698e-08, 
    1.08278e-08, 1.085022e-08, 1.085343e-08, 1.084474e-08, 1.090369e-08, 
    1.088233e-08, 1.093984e-08, 1.09243e-08, 1.094976e-08, 1.093711e-08, 
    1.093525e-08, 1.0919e-08, 1.090888e-08, 1.088331e-08, 1.08625e-08, 
    1.0846e-08, 1.084984e-08, 1.086797e-08, 1.090079e-08, 1.093183e-08, 
    1.092503e-08, 1.094783e-08, 1.088748e-08, 1.091279e-08, 1.090301e-08, 
    1.092851e-08, 1.087263e-08, 1.09202e-08, 1.086046e-08, 1.08657e-08, 
    1.088191e-08, 1.09145e-08, 1.092172e-08, 1.092941e-08, 1.092467e-08, 
    1.090162e-08, 1.089785e-08, 1.088152e-08, 1.087701e-08, 1.086456e-08, 
    1.085426e-08, 1.086367e-08, 1.087356e-08, 1.090163e-08, 1.092693e-08, 
    1.09545e-08, 1.096124e-08, 1.099344e-08, 1.096723e-08, 1.101047e-08, 
    1.09737e-08, 1.103735e-08, 1.092297e-08, 1.097262e-08, 1.088265e-08, 
    1.089235e-08, 1.090988e-08, 1.095009e-08, 1.092839e-08, 1.095377e-08, 
    1.08977e-08, 1.086859e-08, 1.086106e-08, 1.084701e-08, 1.086138e-08, 
    1.086021e-08, 1.087397e-08, 1.086955e-08, 1.090256e-08, 1.088483e-08, 
    1.09352e-08, 1.095357e-08, 1.100545e-08, 1.103724e-08, 1.10696e-08, 
    1.108387e-08, 1.108822e-08, 1.109004e-08 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.200366e-14, 5.213594e-14, 5.211024e-14, 5.221683e-14, 5.215773e-14, 
    5.222749e-14, 5.203051e-14, 5.214117e-14, 5.207055e-14, 5.20156e-14, 
    5.242333e-14, 5.222158e-14, 5.26327e-14, 5.250429e-14, 5.282665e-14, 
    5.26127e-14, 5.286975e-14, 5.282054e-14, 5.296872e-14, 5.292629e-14, 
    5.311549e-14, 5.298829e-14, 5.321352e-14, 5.308516e-14, 5.310523e-14, 
    5.298409e-14, 5.226226e-14, 5.239821e-14, 5.225419e-14, 5.227359e-14, 
    5.226489e-14, 5.215894e-14, 5.210547e-14, 5.199357e-14, 5.20139e-14, 
    5.20961e-14, 5.228231e-14, 5.221917e-14, 5.237833e-14, 5.237474e-14, 
    5.255165e-14, 5.247192e-14, 5.276888e-14, 5.268457e-14, 5.292806e-14, 
    5.286687e-14, 5.292518e-14, 5.290751e-14, 5.292541e-14, 5.283566e-14, 
    5.287412e-14, 5.279512e-14, 5.248685e-14, 5.257752e-14, 5.230685e-14, 
    5.214371e-14, 5.203535e-14, 5.195836e-14, 5.196925e-14, 5.198999e-14, 
    5.209659e-14, 5.219676e-14, 5.227303e-14, 5.232401e-14, 5.237423e-14, 
    5.252597e-14, 5.260631e-14, 5.27859e-14, 5.275355e-14, 5.280837e-14, 
    5.286079e-14, 5.294866e-14, 5.293421e-14, 5.29729e-14, 5.280696e-14, 
    5.291726e-14, 5.273511e-14, 5.278495e-14, 5.238771e-14, 5.223621e-14, 
    5.217162e-14, 5.211518e-14, 5.197762e-14, 5.207262e-14, 5.203518e-14, 
    5.212428e-14, 5.218083e-14, 5.215287e-14, 5.23254e-14, 5.225835e-14, 
    5.261107e-14, 5.245927e-14, 5.285467e-14, 5.276019e-14, 5.287731e-14, 
    5.281757e-14, 5.29199e-14, 5.282781e-14, 5.298731e-14, 5.302199e-14, 
    5.299829e-14, 5.308936e-14, 5.28227e-14, 5.292517e-14, 5.215208e-14, 
    5.215664e-14, 5.21779e-14, 5.208441e-14, 5.20787e-14, 5.199301e-14, 
    5.206928e-14, 5.210173e-14, 5.218412e-14, 5.223281e-14, 5.227908e-14, 
    5.238074e-14, 5.249416e-14, 5.26526e-14, 5.276632e-14, 5.284247e-14, 
    5.279579e-14, 5.2837e-14, 5.279093e-14, 5.276933e-14, 5.300898e-14, 
    5.287447e-14, 5.307626e-14, 5.306511e-14, 5.297381e-14, 5.306637e-14, 
    5.215985e-14, 5.21336e-14, 5.204237e-14, 5.211377e-14, 5.198367e-14, 
    5.205649e-14, 5.209833e-14, 5.225972e-14, 5.229518e-14, 5.232801e-14, 
    5.239286e-14, 5.2476e-14, 5.26217e-14, 5.274834e-14, 5.286384e-14, 
    5.285538e-14, 5.285836e-14, 5.288413e-14, 5.282026e-14, 5.289461e-14, 
    5.290707e-14, 5.287447e-14, 5.306362e-14, 5.300962e-14, 5.306488e-14, 
    5.302972e-14, 5.214213e-14, 5.21863e-14, 5.216243e-14, 5.22073e-14, 
    5.217568e-14, 5.231617e-14, 5.235826e-14, 5.255503e-14, 5.247436e-14, 
    5.260277e-14, 5.248742e-14, 5.250786e-14, 5.260689e-14, 5.249367e-14, 
    5.274133e-14, 5.257342e-14, 5.288513e-14, 5.271761e-14, 5.289562e-14, 
    5.286334e-14, 5.291679e-14, 5.296462e-14, 5.302479e-14, 5.313568e-14, 
    5.311002e-14, 5.320272e-14, 5.225213e-14, 5.230934e-14, 5.230434e-14, 
    5.23642e-14, 5.240845e-14, 5.250434e-14, 5.265792e-14, 5.26002e-14, 
    5.270618e-14, 5.272743e-14, 5.256644e-14, 5.266528e-14, 5.234764e-14, 
    5.239899e-14, 5.236844e-14, 5.225662e-14, 5.261347e-14, 5.243046e-14, 
    5.276819e-14, 5.266923e-14, 5.29578e-14, 5.281435e-14, 5.309589e-14, 
    5.321593e-14, 5.332893e-14, 5.346066e-14, 5.234059e-14, 5.230172e-14, 
    5.237133e-14, 5.246751e-14, 5.255676e-14, 5.267526e-14, 5.26874e-14, 
    5.270957e-14, 5.276703e-14, 5.281529e-14, 5.271655e-14, 5.282739e-14, 
    5.241083e-14, 5.262935e-14, 5.2287e-14, 5.239016e-14, 5.246186e-14, 
    5.243044e-14, 5.259361e-14, 5.263203e-14, 5.278797e-14, 5.27074e-14, 
    5.318629e-14, 5.297468e-14, 5.356095e-14, 5.339743e-14, 5.228813e-14, 
    5.234047e-14, 5.252239e-14, 5.243587e-14, 5.268319e-14, 5.274396e-14, 
    5.279337e-14, 5.285645e-14, 5.286328e-14, 5.290064e-14, 5.283941e-14, 
    5.289823e-14, 5.267552e-14, 5.27751e-14, 5.250164e-14, 5.256825e-14, 
    5.253762e-14, 5.250399e-14, 5.260774e-14, 5.27181e-14, 5.272051e-14, 
    5.275586e-14, 5.285534e-14, 5.268419e-14, 5.321348e-14, 5.288683e-14, 
    5.239751e-14, 5.249813e-14, 5.251255e-14, 5.247358e-14, 5.273787e-14, 
    5.264218e-14, 5.289974e-14, 5.28302e-14, 5.294412e-14, 5.288752e-14, 
    5.287919e-14, 5.280646e-14, 5.276113e-14, 5.264656e-14, 5.255325e-14, 
    5.247924e-14, 5.249646e-14, 5.257775e-14, 5.272486e-14, 5.286388e-14, 
    5.283343e-14, 5.293547e-14, 5.266527e-14, 5.277863e-14, 5.273481e-14, 
    5.284903e-14, 5.259866e-14, 5.281175e-14, 5.254411e-14, 5.256761e-14, 
    5.264028e-14, 5.278628e-14, 5.281863e-14, 5.285307e-14, 5.283183e-14, 
    5.27286e-14, 5.27117e-14, 5.263852e-14, 5.261829e-14, 5.25625e-14, 
    5.251627e-14, 5.25585e-14, 5.260282e-14, 5.272866e-14, 5.284193e-14, 
    5.296529e-14, 5.299548e-14, 5.313928e-14, 5.302217e-14, 5.321529e-14, 
    5.305102e-14, 5.333526e-14, 5.282416e-14, 5.304629e-14, 5.26436e-14, 
    5.268707e-14, 5.276559e-14, 5.294557e-14, 5.284849e-14, 5.296204e-14, 
    5.271104e-14, 5.258053e-14, 5.25468e-14, 5.248373e-14, 5.254824e-14, 
    5.2543e-14, 5.260468e-14, 5.258487e-14, 5.273284e-14, 5.265338e-14, 
    5.287897e-14, 5.296116e-14, 5.319299e-14, 5.333483e-14, 5.347909e-14, 
    5.354268e-14, 5.356204e-14, 5.357012e-14 ;

 POT_F_DENIT =
  2.413656e-36, 2.065401e-35, 1.367197e-35, 7.458777e-35, 2.924233e-35, 
    8.819833e-35, 3.748208e-36, 2.246482e-35, 7.197595e-36, 2.935293e-36, 
    1.796957e-33, 8.037766e-35, 3.922441e-32, 6.007093e-33, 6.052333e-31, 
    2.939911e-32, 1.094422e-30, 5.556852e-31, 4.175555e-30, 2.359349e-30, 
    2.893847e-29, 5.424175e-30, 1.017046e-28, 1.948533e-29, 2.531664e-29, 
    5.128552e-30, 1.5186e-34, 1.229759e-33, 1.339012e-34, 1.812237e-34, 
    1.582295e-34, 2.981927e-35, 1.267358e-35, 2.04289e-36, 2.854736e-36, 
    1.088977e-35, 2.075535e-34, 7.733206e-35, 9.06774e-34, 8.585492e-34, 
    1.206895e-32, 3.712564e-33, 2.708682e-31, 8.236855e-32, 2.416494e-30, 
    1.051322e-30, 2.324528e-30, 1.82943e-30, 2.331775e-30, 6.847458e-31, 
    1.161084e-30, 3.905416e-31, 4.637344e-33, 1.761981e-32, 3.033677e-34, 
    2.342121e-35, 4.05827e-36, 1.140883e-36, 1.366814e-36, 1.926661e-36, 
    1.097471e-35, 5.431533e-35, 1.795261e-34, 3.950291e-34, 8.518304e-34, 
    8.288211e-33, 2.678748e-32, 3.436761e-31, 2.184636e-31, 4.697071e-31, 
    9.671604e-31, 3.190841e-30, 2.625917e-30, 4.41738e-30, 4.603185e-31, 
    2.088884e-30, 1.685259e-31, 3.389846e-31, 1.048926e-33, 1.010662e-34, 
    3.652738e-35, 1.480341e-35, 1.570089e-36, 7.446789e-36, 4.047018e-36, 
    1.712407e-35, 4.221452e-35, 2.705511e-35, 4.035902e-34, 1.42863e-34, 
    2.869719e-32, 3.075397e-33, 8.894096e-31, 2.398156e-31, 1.212633e-30, 
    5.331979e-31, 2.164703e-30, 6.143018e-31, 5.354316e-30, 8.491746e-30, 
    6.198718e-30, 2.057202e-29, 5.724397e-31, 2.324658e-30, 2.671984e-35, 
    2.873639e-35, 4.028986e-35, 9.014748e-36, 8.217192e-36, 2.024267e-36, 
    7.050135e-36, 1.192036e-35, 4.446345e-35, 9.581258e-35, 1.972759e-34, 
    9.40965e-34, 5.171452e-33, 5.218879e-32, 2.613056e-31, 7.518973e-31, 
    3.941118e-31, 6.973537e-31, 3.683514e-31, 2.724792e-31, 7.147453e-30, 
    1.166841e-30, 1.73386e-29, 1.498157e-29, 4.472238e-30, 1.523048e-29, 
    3.024102e-35, 1.988205e-35, 4.550449e-36, 1.44646e-35, 1.73507e-36, 
    5.729078e-36, 1.12904e-35, 1.460426e-34, 2.53197e-34, 4.202358e-34, 
    1.130701e-33, 3.94548e-33, 3.344858e-32, 2.031258e-31, 1.00837e-30, 
    8.979328e-31, 9.353917e-31, 1.33104e-30, 5.534872e-31, 1.535411e-30, 
    1.819247e-30, 1.166494e-30, 1.469084e-29, 7.203947e-30, 1.493503e-29, 
    9.401376e-30, 2.279148e-35, 4.603192e-35, 3.151121e-35, 6.416304e-35, 
    3.891003e-35, 3.504587e-34, 6.685744e-34, 1.269163e-32, 3.850616e-33, 
    2.54377e-32, 4.67595e-33, 6.33306e-33, 2.703684e-32, 5.129652e-33, 
    1.84164e-31, 1.661233e-32, 1.349351e-30, 1.31887e-31, 1.556519e-30, 
    1.001499e-30, 2.074591e-30, 3.953509e-30, 8.809192e-30, 3.754736e-29, 
    2.692728e-29, 8.862534e-29, 1.296324e-34, 3.153121e-34, 2.916695e-34, 
    7.313115e-34, 1.432144e-33, 6.009421e-33, 5.630612e-32, 2.449265e-32, 
    1.119704e-31, 1.512694e-31, 1.497909e-32, 6.257924e-32, 5.680003e-34, 
    1.242106e-33, 7.802933e-34, 1.391165e-34, 2.970523e-32, 1.996976e-33, 
    2.682689e-31, 6.618635e-32, 3.607827e-30, 5.103762e-31, 2.240553e-29, 
    1.049413e-28, 4.315611e-28, 2.151595e-27, 5.097033e-34, 2.801228e-34, 
    8.151042e-34, 3.479038e-33, 1.300711e-32, 7.215027e-32, 8.574919e-32, 
    1.175121e-31, 2.638394e-31, 5.166526e-31, 1.297972e-31, 6.107406e-31, 
    1.487772e-33, 3.735418e-32, 2.231189e-34, 1.086605e-33, 3.196354e-33, 
    1.995071e-33, 2.225378e-32, 3.879716e-32, 3.537037e-31, 1.139286e-31, 
    7.1979e-29, 4.527107e-30, 7.072285e-27, 1.001204e-27, 2.26989e-34, 
    5.086269e-34, 7.850772e-33, 2.164587e-33, 8.075713e-32, 1.909646e-31, 
    3.810726e-31, 9.116114e-31, 1.000794e-30, 1.666826e-30, 7.208881e-31, 
    1.612822e-30, 7.241077e-32, 2.954449e-31, 5.773067e-33, 1.538488e-32, 
    9.818068e-33, 5.978102e-33, 2.731482e-32, 1.326861e-31, 1.371577e-31, 
    2.257592e-31, 9.004322e-31, 8.191729e-32, 1.019036e-28, 1.384652e-30, 
    1.213156e-33, 5.487309e-33, 6.787049e-33, 3.804815e-33, 1.752723e-31, 
    4.491113e-32, 1.646268e-30, 6.348694e-31, 3.001185e-30, 1.393988e-30, 
    1.244232e-30, 4.570806e-31, 2.430007e-31, 4.783712e-32, 1.235653e-32, 
    4.139165e-33, 5.346258e-33, 1.767639e-32, 1.459641e-31, 1.009369e-30, 
    6.642821e-31, 2.670752e-30, 6.253374e-32, 3.104628e-31, 1.679492e-31, 
    8.230366e-31, 2.39545e-32, 4.932957e-31, 1.079973e-32, 1.5238e-32, 
    4.370052e-32, 3.45641e-31, 5.410543e-31, 8.702187e-31, 6.493018e-31, 
    1.538556e-31, 1.211231e-31, 4.260206e-32, 3.183188e-32, 1.413956e-32, 
    7.167403e-33, 1.333833e-32, 2.544929e-32, 1.539362e-31, 7.466343e-31, 
    3.989861e-30, 5.969769e-30, 3.938643e-29, 8.521178e-30, 1.042838e-28, 
    1.24947e-29, 4.677264e-28, 5.850539e-31, 1.171975e-29, 4.582477e-32, 
    8.533778e-32, 2.588349e-31, 3.063866e-30, 8.169875e-31, 3.821891e-30, 
    1.199891e-31, 1.841584e-32, 1.123526e-32, 4.426199e-33, 1.147535e-32, 
    1.062511e-32, 2.613189e-32, 1.959549e-32, 1.632738e-31, 5.273784e-32, 
    1.240751e-30, 3.776026e-30, 7.832231e-29, 4.6458e-28, 2.680098e-27, 
    5.702732e-27, 7.160027e-27, 7.872312e-27 ;

 POT_F_NIT =
  5.750217e-11, 5.781313e-11, 5.775263e-11, 5.800385e-11, 5.786444e-11, 
    5.802901e-11, 5.756515e-11, 5.782544e-11, 5.765922e-11, 5.753012e-11, 
    5.849272e-11, 5.801504e-11, 5.899102e-11, 5.868493e-11, 5.945526e-11, 
    5.894332e-11, 5.955875e-11, 5.944051e-11, 5.979681e-11, 5.969462e-11, 
    6.015131e-11, 5.984398e-11, 6.038875e-11, 6.007787e-11, 6.012642e-11, 
    5.983382e-11, 5.811111e-11, 5.843317e-11, 5.809203e-11, 5.81379e-11, 
    5.811732e-11, 5.786728e-11, 5.774143e-11, 5.747842e-11, 5.752613e-11, 
    5.771934e-11, 5.81585e-11, 5.800927e-11, 5.838576e-11, 5.837725e-11, 
    5.879765e-11, 5.860792e-11, 5.931663e-11, 5.911481e-11, 5.969888e-11, 
    5.955173e-11, 5.969195e-11, 5.964942e-11, 5.969249e-11, 5.947676e-11, 
    5.956913e-11, 5.937948e-11, 5.864348e-11, 5.885935e-11, 5.821654e-11, 
    5.783151e-11, 5.757652e-11, 5.739587e-11, 5.742138e-11, 5.747004e-11, 
    5.772046e-11, 5.795639e-11, 5.813648e-11, 5.825707e-11, 5.837602e-11, 
    5.873661e-11, 5.892799e-11, 5.935744e-11, 5.927987e-11, 5.941133e-11, 
    5.95371e-11, 5.974848e-11, 5.971366e-11, 5.980686e-11, 5.940787e-11, 
    5.967288e-11, 5.923566e-11, 5.935508e-11, 5.840826e-11, 5.804954e-11, 
    5.789725e-11, 5.77642e-11, 5.7441e-11, 5.766409e-11, 5.757609e-11, 
    5.778556e-11, 5.791883e-11, 5.78529e-11, 5.826037e-11, 5.810179e-11, 
    5.893933e-11, 5.85779e-11, 5.952243e-11, 5.929578e-11, 5.95768e-11, 
    5.943333e-11, 5.967924e-11, 5.94579e-11, 5.984158e-11, 5.992525e-11, 
    5.986805e-11, 6.008793e-11, 5.944561e-11, 5.969188e-11, 5.785108e-11, 
    5.786183e-11, 5.791192e-11, 5.769182e-11, 5.767837e-11, 5.747708e-11, 
    5.765617e-11, 5.773251e-11, 5.792656e-11, 5.804145e-11, 5.815077e-11, 
    5.839148e-11, 5.866082e-11, 5.903844e-11, 5.931045e-11, 5.949308e-11, 
    5.938107e-11, 5.947995e-11, 5.936941e-11, 5.931762e-11, 5.989387e-11, 
    5.956997e-11, 6.005627e-11, 6.002932e-11, 5.980904e-11, 6.003234e-11, 
    5.786937e-11, 5.780751e-11, 5.759297e-11, 5.776083e-11, 5.745516e-11, 
    5.762614e-11, 5.772455e-11, 5.810506e-11, 5.818885e-11, 5.826654e-11, 
    5.842018e-11, 5.861759e-11, 5.896465e-11, 5.926738e-11, 5.954441e-11, 
    5.952409e-11, 5.953123e-11, 5.959317e-11, 5.943977e-11, 5.961836e-11, 
    5.964834e-11, 5.956993e-11, 6.00257e-11, 5.989533e-11, 6.002873e-11, 
    5.994383e-11, 5.782761e-11, 5.793171e-11, 5.787544e-11, 5.798126e-11, 
    5.790668e-11, 5.823857e-11, 5.833824e-11, 5.880572e-11, 5.86137e-11, 
    5.891949e-11, 5.864472e-11, 5.869336e-11, 5.89294e-11, 5.865956e-11, 
    5.925063e-11, 5.884954e-11, 5.959556e-11, 5.919391e-11, 5.962077e-11, 
    5.954317e-11, 5.967168e-11, 5.978686e-11, 5.993194e-11, 6.020002e-11, 
    6.013789e-11, 6.036242e-11, 5.808708e-11, 5.822239e-11, 5.821049e-11, 
    5.835225e-11, 5.845719e-11, 5.868497e-11, 5.905113e-11, 5.891332e-11, 
    5.916644e-11, 5.92173e-11, 5.883279e-11, 5.906871e-11, 5.8313e-11, 
    5.843476e-11, 5.836226e-11, 5.809767e-11, 5.894497e-11, 5.850941e-11, 
    5.931489e-11, 5.907807e-11, 5.977041e-11, 5.94256e-11, 6.01037e-11, 
    6.039458e-11, 6.066907e-11, 6.099039e-11, 5.829632e-11, 5.82043e-11, 
    5.836913e-11, 5.859747e-11, 5.880978e-11, 5.909255e-11, 5.912153e-11, 
    5.917457e-11, 5.93121e-11, 5.942784e-11, 5.91913e-11, 5.945686e-11, 
    5.846295e-11, 5.898286e-11, 5.816944e-11, 5.841379e-11, 5.858394e-11, 
    5.85093e-11, 5.889752e-11, 5.898917e-11, 5.93623e-11, 5.916929e-11, 
    6.032268e-11, 5.981113e-11, 6.123567e-11, 6.083601e-11, 5.817216e-11, 
    5.8296e-11, 5.872794e-11, 5.852224e-11, 5.911145e-11, 5.925688e-11, 
    5.937525e-11, 5.952668e-11, 5.954305e-11, 5.963287e-11, 5.94857e-11, 
    5.962705e-11, 5.90931e-11, 5.933144e-11, 5.867847e-11, 5.883707e-11, 
    5.876409e-11, 5.868406e-11, 5.893119e-11, 5.919495e-11, 5.920064e-11, 
    5.928532e-11, 5.952417e-11, 5.911376e-11, 6.038874e-11, 5.959979e-11, 
    5.843118e-11, 5.867026e-11, 5.87045e-11, 5.86118e-11, 5.924228e-11, 
    5.901347e-11, 5.963068e-11, 5.946359e-11, 5.973748e-11, 5.96013e-11, 
    5.958126e-11, 5.94066e-11, 5.929796e-11, 5.902391e-11, 5.880135e-11, 
    5.862519e-11, 5.866613e-11, 5.885972e-11, 5.921111e-11, 5.954445e-11, 
    5.947134e-11, 5.971658e-11, 5.906854e-11, 5.933986e-11, 5.92349e-11, 
    5.950873e-11, 5.890963e-11, 5.941956e-11, 5.877958e-11, 5.883557e-11, 
    5.900892e-11, 5.935832e-11, 5.943581e-11, 5.951852e-11, 5.946747e-11, 
    5.922009e-11, 5.917961e-11, 5.900468e-11, 5.89564e-11, 5.882334e-11, 
    5.871324e-11, 5.881381e-11, 5.891948e-11, 5.922017e-11, 5.949172e-11, 
    5.978843e-11, 5.986117e-11, 6.020878e-11, 5.992568e-11, 6.039312e-11, 
    5.999549e-11, 6.068461e-11, 5.944924e-11, 5.9984e-11, 5.901683e-11, 
    5.912069e-11, 5.93087e-11, 5.974105e-11, 5.95075e-11, 5.978069e-11, 
    5.917803e-11, 5.886639e-11, 5.878593e-11, 5.863588e-11, 5.878936e-11, 
    5.877687e-11, 5.892389e-11, 5.887662e-11, 5.923016e-11, 5.904013e-11, 
    5.958068e-11, 5.977849e-11, 6.03388e-11, 6.068343e-11, 6.103525e-11, 
    6.119084e-11, 6.123824e-11, 6.125805e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005836714, 0.0005836741, 0.0005836736, 0.0005836757, 0.0005836746, 
    0.000583676, 0.000583672, 0.0005836742, 0.0005836728, 0.0005836717, 
    0.0005836799, 0.0005836759, 0.0005836804, 0.0005836817, 0.0005836844, 
    0.0005836799, 0.0005836854, 0.0005836844, 0.0005836874, 0.0005836866, 
    0.0005836905, 0.0005836879, 0.0005836926, 0.0005836899, 0.0005836902, 
    0.0005836878, 0.0005836767, 0.0005836794, 0.0005836766, 0.000583677, 
    0.0005836768, 0.0005836746, 0.0005836735, 0.0005836712, 0.0005836716, 
    0.0005836733, 0.0005836771, 0.0005836759, 0.0005836792, 0.0005836791, 
    0.0005836827, 0.0005836811, 0.0005836833, 0.0005836816, 0.0005836866, 
    0.0005836854, 0.0005836866, 0.0005836862, 0.0005836866, 0.0005836847, 
    0.0005836855, 0.0005836838, 0.0005836814, 0.0005836793, 0.0005836777, 
    0.0005836742, 0.0005836721, 0.0005836705, 0.0005836707, 0.0005836711, 
    0.0005836733, 0.0005836754, 0.000583677, 0.000583678, 0.0005836791, 
    0.0005836821, 0.0005836798, 0.0005836836, 0.000583683, 0.0005836841, 
    0.0005836852, 0.000583687, 0.0005836867, 0.0005836876, 0.0005836841, 
    0.0005836863, 0.0005836826, 0.0005836836, 0.0005836792, 0.0005836762, 
    0.0005836748, 0.0005836737, 0.0005836709, 0.0005836728, 0.000583672, 
    0.0005836739, 0.000583675, 0.0005836745, 0.0005836781, 0.0005836767, 
    0.0005836799, 0.0005836808, 0.0005836851, 0.0005836831, 0.0005836856, 
    0.0005836843, 0.0005836864, 0.0005836845, 0.0005836879, 0.0005836886, 
    0.0005836881, 0.00058369, 0.0005836844, 0.0005836865, 0.0005836745, 
    0.0005836746, 0.000583675, 0.0005836731, 0.000583673, 0.0005836712, 
    0.0005836728, 0.0005836734, 0.0005836752, 0.0005836762, 0.0005836771, 
    0.0005836792, 0.0005836815, 0.0005836808, 0.0005836833, 0.0005836848, 
    0.0005836838, 0.0005836847, 0.0005836838, 0.0005836833, 0.0005836883, 
    0.0005836855, 0.0005836897, 0.0005836895, 0.0005836876, 0.0005836895, 
    0.0005836746, 0.0005836741, 0.0005836722, 0.0005836737, 0.000583671, 
    0.0005836725, 0.0005836733, 0.0005836767, 0.0005836774, 0.0005836781, 
    0.0005836795, 0.0005836812, 0.0005836802, 0.0005836828, 0.0005836853, 
    0.0005836851, 0.0005836852, 0.0005836857, 0.0005836844, 0.0005836859, 
    0.0005836862, 0.0005836855, 0.0005836895, 0.0005836883, 0.0005836895, 
    0.0005836887, 0.0005836743, 0.0005836752, 0.0005836747, 0.0005836756, 
    0.0005836749, 0.0005836778, 0.0005836787, 0.0005836827, 0.0005836811, 
    0.0005836798, 0.0005836814, 0.0005836818, 0.0005836798, 0.0005836815, 
    0.0005836827, 0.0005836791, 0.0005836857, 0.0005836821, 0.0005836859, 
    0.0005836853, 0.0005836864, 0.0005836874, 0.0005836887, 0.0005836909, 
    0.0005836904, 0.0005836923, 0.0005836766, 0.0005836777, 0.0005836776, 
    0.0005836788, 0.0005836798, 0.0005836817, 0.000583681, 0.0005836798, 
    0.000583682, 0.0005836824, 0.0005836791, 0.0005836811, 0.0005836785, 
    0.0005836795, 0.0005836789, 0.0005836766, 0.00058368, 0.0005836802, 
    0.0005836833, 0.0005836812, 0.0005836872, 0.0005836842, 0.0005836901, 
    0.0005836926, 0.000583695, 0.0005836978, 0.0005836784, 0.0005836776, 
    0.000583679, 0.0005836809, 0.0005836789, 0.0005836813, 0.0005836816, 
    0.000583682, 0.0005836833, 0.0005836842, 0.0005836822, 0.0005836845, 
    0.0005836796, 0.0005836803, 0.0005836773, 0.0005836793, 0.0005836808, 
    0.0005836802, 0.0005836796, 0.0005836805, 0.0005836837, 0.000583682, 
    0.0005836919, 0.0005836875, 0.0005836999, 0.0005836964, 0.0005836773, 
    0.0005836784, 0.0005836821, 0.0005836803, 0.0005836815, 0.0005836828, 
    0.0005836838, 0.0005836851, 0.0005836853, 0.0005836861, 0.0005836848, 
    0.000583686, 0.0005836813, 0.0005836834, 0.0005836817, 0.0005836791, 
    0.0005836824, 0.0005836817, 0.0005836799, 0.0005836822, 0.0005836823, 
    0.000583683, 0.0005836849, 0.0005836815, 0.0005836924, 0.0005836856, 
    0.0005836795, 0.0005836816, 0.0005836819, 0.0005836811, 0.0005836826, 
    0.0005836806, 0.000583686, 0.0005836846, 0.000583687, 0.0005836858, 
    0.0005836856, 0.0005836841, 0.0005836831, 0.0005836808, 0.0005836827, 
    0.0005836812, 0.0005836816, 0.0005836793, 0.0005836823, 0.0005836852, 
    0.0005836846, 0.0005836867, 0.0005836812, 0.0005836835, 0.0005836826, 
    0.0005836849, 0.0005836798, 0.000583684, 0.0005836826, 0.0005836791, 
    0.0005836806, 0.0005836836, 0.0005836844, 0.000583685, 0.0005836846, 
    0.0005836824, 0.0005836821, 0.0005836806, 0.0005836802, 0.000583679, 
    0.000583682, 0.0005836789, 0.0005836798, 0.0005836824, 0.0005836848, 
    0.0005836874, 0.000583688, 0.0005836909, 0.0005836885, 0.0005836924, 
    0.000583689, 0.000583695, 0.0005836844, 0.000583689, 0.0005836807, 
    0.0005836816, 0.0005836832, 0.0005836869, 0.0005836849, 0.0005836873, 
    0.0005836821, 0.0005836793, 0.0005836826, 0.0005836813, 0.0005836827, 
    0.0005836826, 0.0005836799, 0.0005836795, 0.0005836826, 0.0005836809, 
    0.0005836856, 0.0005836873, 0.0005836921, 0.0005836951, 0.0005836982, 
    0.0005836996, 0.0005837, 0.0005837001 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_NODYNLNDUSE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_R =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.18217, 81.18126, 81.18143, 81.18071, 81.18111, 81.18064, 81.18198, 
    81.18123, 81.1817, 81.18208, 81.17934, 81.18068, 81.17746, 81.17873, 
    81.17612, 81.17761, 81.17582, 81.17615, 81.17511, 81.17541, 81.17413, 
    81.17498, 81.17343, 81.17432, 81.17419, 81.17501, 81.18039, 81.17951, 
    81.18044, 81.18032, 81.18037, 81.18111, 81.18148, 81.18222, 81.18208, 
    81.18153, 81.18026, 81.18068, 81.17959, 81.17961, 81.17841, 81.17895, 
    81.17651, 81.17708, 81.17539, 81.17582, 81.17542, 81.17554, 81.17542, 
    81.17604, 81.17577, 81.17632, 81.17885, 81.17783, 81.18009, 81.18124, 
    81.18195, 81.18246, 81.18239, 81.18225, 81.18153, 81.18083, 81.18031, 
    81.17996, 81.17962, 81.17862, 81.17764, 81.1764, 81.17661, 81.17624, 
    81.17587, 81.17525, 81.17535, 81.17509, 81.17624, 81.17548, 81.17673, 
    81.17639, 81.17959, 81.18056, 81.18104, 81.1814, 81.18233, 81.18169, 
    81.18195, 81.18133, 81.18095, 81.18113, 81.17995, 81.18041, 81.17761, 
    81.17905, 81.17591, 81.17656, 81.17575, 81.17616, 81.17546, 81.17609, 
    81.17499, 81.17476, 81.17492, 81.17428, 81.17612, 81.17542, 81.18114, 
    81.18111, 81.18096, 81.18162, 81.18165, 81.18223, 81.18171, 81.1815, 
    81.18092, 81.18059, 81.18027, 81.17958, 81.17881, 81.17731, 81.17652, 
    81.17599, 81.17631, 81.17603, 81.17635, 81.17649, 81.17485, 81.17577, 
    81.17437, 81.17445, 81.17509, 81.17444, 81.18109, 81.18127, 81.18189, 
    81.1814, 81.18229, 81.1818, 81.18153, 81.18042, 81.18016, 81.17994, 
    81.17949, 81.17892, 81.17753, 81.17665, 81.17584, 81.1759, 81.17588, 
    81.1757, 81.17615, 81.17563, 81.17555, 81.17577, 81.17445, 81.17483, 
    81.17445, 81.17469, 81.18121, 81.18091, 81.18107, 81.18077, 81.18098, 
    81.18004, 81.17975, 81.1784, 81.17894, 81.17766, 81.17884, 81.17871, 
    81.17766, 81.17879, 81.17671, 81.17788, 81.1757, 81.17689, 81.17562, 
    81.17584, 81.17548, 81.17515, 81.17473, 81.17397, 81.17414, 81.17349, 
    81.18046, 81.18008, 81.1801, 81.17969, 81.17939, 81.17873, 81.17727, 
    81.17767, 81.17693, 81.17679, 81.17789, 81.17722, 81.17981, 81.17947, 
    81.17966, 81.18044, 81.17759, 81.17925, 81.17651, 81.17719, 81.17519, 
    81.1762, 81.17424, 81.17343, 81.17261, 81.17172, 81.17986, 81.18011, 
    81.17963, 81.179, 81.17797, 81.17715, 81.17706, 81.17691, 81.17651, 
    81.17618, 81.17688, 81.17609, 81.17942, 81.17747, 81.18022, 81.17953, 
    81.17903, 81.17924, 81.1777, 81.17744, 81.17638, 81.17692, 81.17365, 
    81.17509, 81.171, 81.17216, 81.18021, 81.17985, 81.17861, 81.1792, 
    81.17709, 81.17667, 81.17632, 81.1759, 81.17584, 81.17559, 81.17601, 
    81.17561, 81.17715, 81.17646, 81.17874, 81.17789, 81.17849, 81.17873, 
    81.17761, 81.17687, 81.17683, 81.1766, 81.17597, 81.17709, 81.17349, 
    81.17575, 81.17946, 81.17879, 81.17867, 81.17893, 81.17672, 81.17738, 
    81.1756, 81.17607, 81.17529, 81.17567, 81.17574, 81.17624, 81.17655, 
    81.17735, 81.1784, 81.17889, 81.17878, 81.17783, 81.17682, 81.17585, 
    81.17606, 81.17535, 81.17722, 81.17645, 81.17675, 81.17595, 81.17768, 
    81.17626, 81.17844, 81.17789, 81.17739, 81.1764, 81.17616, 81.17593, 
    81.17606, 81.17679, 81.1769, 81.1774, 81.17754, 81.17792, 81.17864, 
    81.17795, 81.17766, 81.17678, 81.176, 81.17515, 81.17493, 81.17397, 
    81.17478, 81.17348, 81.17463, 81.17262, 81.17616, 81.17462, 81.17736, 
    81.17706, 81.17654, 81.1753, 81.17595, 81.17518, 81.1769, 81.17782, 
    81.17843, 81.17886, 81.17842, 81.17846, 81.17763, 81.17776, 81.17675, 
    81.17729, 81.17574, 81.17519, 81.17357, 81.17259, 81.17156, 81.17112, 
    81.17098, 81.17092 ;

 RH2M_R =
  81.18217, 81.18126, 81.18143, 81.18071, 81.18111, 81.18064, 81.18198, 
    81.18123, 81.1817, 81.18208, 81.17934, 81.18068, 81.17746, 81.17873, 
    81.17612, 81.17761, 81.17582, 81.17615, 81.17511, 81.17541, 81.17413, 
    81.17498, 81.17343, 81.17432, 81.17419, 81.17501, 81.18039, 81.17951, 
    81.18044, 81.18032, 81.18037, 81.18111, 81.18148, 81.18222, 81.18208, 
    81.18153, 81.18026, 81.18068, 81.17959, 81.17961, 81.17841, 81.17895, 
    81.17651, 81.17708, 81.17539, 81.17582, 81.17542, 81.17554, 81.17542, 
    81.17604, 81.17577, 81.17632, 81.17885, 81.17783, 81.18009, 81.18124, 
    81.18195, 81.18246, 81.18239, 81.18225, 81.18153, 81.18083, 81.18031, 
    81.17996, 81.17962, 81.17862, 81.17764, 81.1764, 81.17661, 81.17624, 
    81.17587, 81.17525, 81.17535, 81.17509, 81.17624, 81.17548, 81.17673, 
    81.17639, 81.17959, 81.18056, 81.18104, 81.1814, 81.18233, 81.18169, 
    81.18195, 81.18133, 81.18095, 81.18113, 81.17995, 81.18041, 81.17761, 
    81.17905, 81.17591, 81.17656, 81.17575, 81.17616, 81.17546, 81.17609, 
    81.17499, 81.17476, 81.17492, 81.17428, 81.17612, 81.17542, 81.18114, 
    81.18111, 81.18096, 81.18162, 81.18165, 81.18223, 81.18171, 81.1815, 
    81.18092, 81.18059, 81.18027, 81.17958, 81.17881, 81.17731, 81.17652, 
    81.17599, 81.17631, 81.17603, 81.17635, 81.17649, 81.17485, 81.17577, 
    81.17437, 81.17445, 81.17509, 81.17444, 81.18109, 81.18127, 81.18189, 
    81.1814, 81.18229, 81.1818, 81.18153, 81.18042, 81.18016, 81.17994, 
    81.17949, 81.17892, 81.17753, 81.17665, 81.17584, 81.1759, 81.17588, 
    81.1757, 81.17615, 81.17563, 81.17555, 81.17577, 81.17445, 81.17483, 
    81.17445, 81.17469, 81.18121, 81.18091, 81.18107, 81.18077, 81.18098, 
    81.18004, 81.17975, 81.1784, 81.17894, 81.17766, 81.17884, 81.17871, 
    81.17766, 81.17879, 81.17671, 81.17788, 81.1757, 81.17689, 81.17562, 
    81.17584, 81.17548, 81.17515, 81.17473, 81.17397, 81.17414, 81.17349, 
    81.18046, 81.18008, 81.1801, 81.17969, 81.17939, 81.17873, 81.17727, 
    81.17767, 81.17693, 81.17679, 81.17789, 81.17722, 81.17981, 81.17947, 
    81.17966, 81.18044, 81.17759, 81.17925, 81.17651, 81.17719, 81.17519, 
    81.1762, 81.17424, 81.17343, 81.17261, 81.17172, 81.17986, 81.18011, 
    81.17963, 81.179, 81.17797, 81.17715, 81.17706, 81.17691, 81.17651, 
    81.17618, 81.17688, 81.17609, 81.17942, 81.17747, 81.18022, 81.17953, 
    81.17903, 81.17924, 81.1777, 81.17744, 81.17638, 81.17692, 81.17365, 
    81.17509, 81.171, 81.17216, 81.18021, 81.17985, 81.17861, 81.1792, 
    81.17709, 81.17667, 81.17632, 81.1759, 81.17584, 81.17559, 81.17601, 
    81.17561, 81.17715, 81.17646, 81.17874, 81.17789, 81.17849, 81.17873, 
    81.17761, 81.17687, 81.17683, 81.1766, 81.17597, 81.17709, 81.17349, 
    81.17575, 81.17946, 81.17879, 81.17867, 81.17893, 81.17672, 81.17738, 
    81.1756, 81.17607, 81.17529, 81.17567, 81.17574, 81.17624, 81.17655, 
    81.17735, 81.1784, 81.17889, 81.17878, 81.17783, 81.17682, 81.17585, 
    81.17606, 81.17535, 81.17722, 81.17645, 81.17675, 81.17595, 81.17768, 
    81.17626, 81.17844, 81.17789, 81.17739, 81.1764, 81.17616, 81.17593, 
    81.17606, 81.17679, 81.1769, 81.1774, 81.17754, 81.17792, 81.17864, 
    81.17795, 81.17766, 81.17678, 81.176, 81.17515, 81.17493, 81.17397, 
    81.17478, 81.17348, 81.17463, 81.17262, 81.17616, 81.17462, 81.17736, 
    81.17706, 81.17654, 81.1753, 81.17595, 81.17518, 81.1769, 81.17782, 
    81.17843, 81.17886, 81.17842, 81.17846, 81.17763, 81.17776, 81.17675, 
    81.17729, 81.17574, 81.17519, 81.17357, 81.17259, 81.17156, 81.17112, 
    81.17098, 81.17092 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RSCANOPY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0005333438, 0.000534749, 0.0005344758, 0.0005356089, 0.0005349804, 
    0.0005357221, 0.0005336285, 0.0005348044, 0.0005340537, 0.00053347, 
    0.0005378062, 0.000535659, 0.0005400364, 0.0005386675, 0.0005421054, 
    0.0005398232, 0.0005425653, 0.0005420396, 0.000543622, 0.0005431686, 
    0.0005451916, 0.0005438311, 0.0005462401, 0.0005448668, 0.0005450814, 
    0.0005437859, 0.0005360918, 0.0005375394, 0.0005360059, 0.0005362123, 
    0.0005361197, 0.0005349931, 0.0005344251, 0.000533236, 0.0005334519, 
    0.0005343253, 0.0005363048, 0.0005356329, 0.000537326, 0.0005372879, 
    0.0005391719, 0.0005383225, 0.0005414882, 0.0005405886, 0.0005431875, 
    0.0005425339, 0.0005431567, 0.0005429678, 0.000543159, 0.0005422006, 
    0.0005426111, 0.0005417677, 0.0005384822, 0.0005394482, 0.000536566, 
    0.0005348317, 0.0005336798, 0.0005328622, 0.0005329777, 0.000533198, 
    0.0005343303, 0.0005353946, 0.0005362056, 0.0005367479, 0.0005372822, 
    0.0005388988, 0.0005397546, 0.0005416698, 0.0005413244, 0.0005419096, 
    0.0005424689, 0.0005434075, 0.000543253, 0.0005436663, 0.000541894, 
    0.0005430719, 0.0005411271, 0.0005416591, 0.0005374274, 0.0005358144, 
    0.0005351282, 0.0005345278, 0.0005330665, 0.0005340756, 0.0005336778, 
    0.0005346242, 0.0005352253, 0.0005349279, 0.0005367626, 0.0005360493, 
    0.0005398052, 0.0005381878, 0.0005424037, 0.0005413952, 0.0005426452, 
    0.0005420074, 0.0005431001, 0.0005421166, 0.0005438201, 0.000544191, 
    0.0005439374, 0.000544911, 0.0005420618, 0.0005431561, 0.0005349199, 
    0.0005349684, 0.0005351942, 0.0005342009, 0.0005341401, 0.0005332297, 
    0.0005340397, 0.0005343846, 0.0005352601, 0.0005357777, 0.0005362697, 
    0.0005373515, 0.0005385593, 0.0005402477, 0.0005414605, 0.0005422731, 
    0.0005417748, 0.0005422147, 0.0005417228, 0.0005414922, 0.0005440518, 
    0.0005426147, 0.0005447709, 0.0005446516, 0.0005436757, 0.0005446649, 
    0.0005350023, 0.0005347232, 0.000533754, 0.0005345124, 0.0005331304, 
    0.0005339039, 0.0005343485, 0.000536064, 0.0005364409, 0.0005367903, 
    0.0005374803, 0.0005383655, 0.0005399181, 0.0005412686, 0.0005425012, 
    0.0005424108, 0.0005424426, 0.0005427178, 0.0005420358, 0.0005428296, 
    0.0005429627, 0.0005426144, 0.0005446355, 0.0005440582, 0.0005446489, 
    0.0005442729, 0.0005348139, 0.0005352833, 0.0005350295, 0.0005355066, 
    0.0005351703, 0.0005366646, 0.0005371125, 0.0005392078, 0.000538348, 
    0.0005397164, 0.000538487, 0.0005387049, 0.0005397606, 0.0005385533, 
    0.0005411939, 0.0005394035, 0.0005427284, 0.000540941, 0.0005428403, 
    0.0005424955, 0.0005430662, 0.0005435773, 0.0005442202, 0.0005454063, 
    0.0005451316, 0.0005461234, 0.0005359832, 0.0005365919, 0.0005365384, 
    0.0005371754, 0.0005376464, 0.0005386674, 0.0005403043, 0.0005396888, 
    0.0005408186, 0.0005410454, 0.0005393287, 0.0005403826, 0.0005369988, 
    0.0005375454, 0.00053722, 0.0005360303, 0.00053983, 0.0005378802, 
    0.0005414799, 0.0005404241, 0.0005435043, 0.0005419726, 0.0005449803, 
    0.0005462653, 0.0005474747, 0.000548887, 0.0005369242, 0.0005365104, 
    0.0005372511, 0.0005382754, 0.0005392259, 0.0005404891, 0.0005406184, 
    0.0005408548, 0.0005414676, 0.0005419828, 0.0005409294, 0.0005421118, 
    0.000537672, 0.0005399992, 0.0005363532, 0.0005374512, 0.0005382143, 
    0.0005378797, 0.0005396177, 0.0005400272, 0.0005416907, 0.0005408309, 
    0.0005459479, 0.0005436847, 0.0005499624, 0.0005482089, 0.0005363658, 
    0.0005369225, 0.0005388596, 0.0005379381, 0.0005405733, 0.0005412218, 
    0.0005417488, 0.0005424223, 0.000542495, 0.000542894, 0.00054224, 
    0.0005428682, 0.0005404913, 0.0005415535, 0.0005386378, 0.0005393475, 
    0.000539021, 0.0005386627, 0.0005397681, 0.0005409453, 0.0005409706, 
    0.0005413479, 0.0005424107, 0.000540583, 0.0005462393, 0.0005427466, 
    0.0005375296, 0.0005386014, 0.0005387546, 0.0005383394, 0.0005411566, 
    0.000540136, 0.0005428843, 0.0005421417, 0.0005433583, 0.0005427537, 
    0.0005426647, 0.0005418881, 0.0005414044, 0.0005401823, 0.0005391877, 
    0.000538399, 0.0005385823, 0.0005394486, 0.0005410172, 0.0005425008, 
    0.0005421758, 0.0005432651, 0.0005403812, 0.0005415906, 0.000541123, 
    0.0005423418, 0.0005396722, 0.000541946, 0.0005390906, 0.000539341, 
    0.0005401156, 0.0005416733, 0.000542018, 0.0005423859, 0.0005421588, 
    0.0005410575, 0.000540877, 0.0005400964, 0.0005398807, 0.000539286, 
    0.0005387933, 0.0005392433, 0.0005397157, 0.0005410576, 0.0005422664, 
    0.0005435839, 0.0005439064, 0.0005454447, 0.0005441921, 0.0005462585, 
    0.0005445012, 0.0005475428, 0.0005420779, 0.000544451, 0.0005401509, 
    0.0005406143, 0.0005414523, 0.0005433741, 0.0005423368, 0.0005435499, 
    0.0005408699, 0.0005394786, 0.0005391186, 0.0005384469, 0.0005391338, 
    0.000539078, 0.0005397354, 0.0005395241, 0.000541102, 0.0005402545, 
    0.0005426616, 0.0005435398, 0.0005460188, 0.0005475376, 0.0005490835, 
    0.0005497657, 0.0005499733, 0.0005500601 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.610009e-14, 3.619188e-14, 3.617406e-14, 3.624802e-14, 3.620701e-14, 
    3.625542e-14, 3.611872e-14, 3.619551e-14, 3.614651e-14, 3.610838e-14, 
    3.639132e-14, 3.625132e-14, 3.653662e-14, 3.644751e-14, 3.667121e-14, 
    3.652274e-14, 3.670112e-14, 3.666697e-14, 3.67698e-14, 3.674036e-14, 
    3.687166e-14, 3.678338e-14, 3.693968e-14, 3.685061e-14, 3.686453e-14, 
    3.678046e-14, 3.627955e-14, 3.63739e-14, 3.627395e-14, 3.628741e-14, 
    3.628138e-14, 3.620785e-14, 3.617075e-14, 3.609309e-14, 3.61072e-14, 
    3.616424e-14, 3.629346e-14, 3.624965e-14, 3.63601e-14, 3.635761e-14, 
    3.648037e-14, 3.642505e-14, 3.663112e-14, 3.657262e-14, 3.674159e-14, 
    3.669912e-14, 3.673959e-14, 3.672732e-14, 3.673975e-14, 3.667746e-14, 
    3.670415e-14, 3.664933e-14, 3.64354e-14, 3.649833e-14, 3.631049e-14, 
    3.619729e-14, 3.612209e-14, 3.606866e-14, 3.607621e-14, 3.609061e-14, 
    3.616458e-14, 3.623409e-14, 3.628702e-14, 3.63224e-14, 3.635725e-14, 
    3.646255e-14, 3.65183e-14, 3.664293e-14, 3.662048e-14, 3.665853e-14, 
    3.66949e-14, 3.675588e-14, 3.674585e-14, 3.67727e-14, 3.665755e-14, 
    3.673409e-14, 3.660769e-14, 3.664228e-14, 3.636661e-14, 3.626147e-14, 
    3.621665e-14, 3.617748e-14, 3.608202e-14, 3.614795e-14, 3.612196e-14, 
    3.618379e-14, 3.622304e-14, 3.620364e-14, 3.632337e-14, 3.627684e-14, 
    3.65216e-14, 3.641627e-14, 3.669066e-14, 3.662509e-14, 3.670637e-14, 
    3.666491e-14, 3.673592e-14, 3.667202e-14, 3.67827e-14, 3.680677e-14, 
    3.679032e-14, 3.685352e-14, 3.666847e-14, 3.673958e-14, 3.620309e-14, 
    3.620625e-14, 3.622101e-14, 3.615613e-14, 3.615217e-14, 3.60927e-14, 
    3.614563e-14, 3.616814e-14, 3.622533e-14, 3.625911e-14, 3.629122e-14, 
    3.636177e-14, 3.644048e-14, 3.655043e-14, 3.662934e-14, 3.668219e-14, 
    3.66498e-14, 3.66784e-14, 3.664642e-14, 3.663143e-14, 3.679774e-14, 
    3.670439e-14, 3.684443e-14, 3.683669e-14, 3.677334e-14, 3.683756e-14, 
    3.620848e-14, 3.619026e-14, 3.612695e-14, 3.61765e-14, 3.608622e-14, 
    3.613676e-14, 3.616579e-14, 3.627778e-14, 3.63024e-14, 3.632518e-14, 
    3.637018e-14, 3.642788e-14, 3.652898e-14, 3.661687e-14, 3.669702e-14, 
    3.669115e-14, 3.669322e-14, 3.67111e-14, 3.666678e-14, 3.671837e-14, 
    3.672702e-14, 3.67044e-14, 3.683566e-14, 3.679818e-14, 3.683653e-14, 
    3.681213e-14, 3.619619e-14, 3.622684e-14, 3.621028e-14, 3.624141e-14, 
    3.621947e-14, 3.631696e-14, 3.634617e-14, 3.648272e-14, 3.642673e-14, 
    3.651585e-14, 3.64358e-14, 3.644998e-14, 3.651871e-14, 3.644014e-14, 
    3.6612e-14, 3.649548e-14, 3.671179e-14, 3.659555e-14, 3.671907e-14, 
    3.669667e-14, 3.673377e-14, 3.676696e-14, 3.680871e-14, 3.688567e-14, 
    3.686786e-14, 3.693218e-14, 3.627252e-14, 3.631222e-14, 3.630875e-14, 
    3.635029e-14, 3.6381e-14, 3.644754e-14, 3.655412e-14, 3.651407e-14, 
    3.658761e-14, 3.660236e-14, 3.649064e-14, 3.655923e-14, 3.63388e-14, 
    3.637443e-14, 3.635323e-14, 3.627564e-14, 3.652327e-14, 3.639627e-14, 
    3.663064e-14, 3.656197e-14, 3.676222e-14, 3.666268e-14, 3.685805e-14, 
    3.694136e-14, 3.701977e-14, 3.711119e-14, 3.633391e-14, 3.630694e-14, 
    3.635524e-14, 3.642198e-14, 3.648392e-14, 3.656615e-14, 3.657458e-14, 
    3.658996e-14, 3.662983e-14, 3.666333e-14, 3.659481e-14, 3.667173e-14, 
    3.638265e-14, 3.65343e-14, 3.629672e-14, 3.63683e-14, 3.641806e-14, 
    3.639626e-14, 3.65095e-14, 3.653615e-14, 3.664437e-14, 3.658846e-14, 
    3.692078e-14, 3.677394e-14, 3.718078e-14, 3.70673e-14, 3.62975e-14, 
    3.633382e-14, 3.646007e-14, 3.640003e-14, 3.657165e-14, 3.661383e-14, 
    3.664812e-14, 3.669189e-14, 3.669663e-14, 3.672256e-14, 3.668007e-14, 
    3.672089e-14, 3.656633e-14, 3.663544e-14, 3.644567e-14, 3.649189e-14, 
    3.647064e-14, 3.64473e-14, 3.651929e-14, 3.659588e-14, 3.659755e-14, 
    3.662209e-14, 3.669112e-14, 3.657235e-14, 3.693965e-14, 3.671297e-14, 
    3.637341e-14, 3.644323e-14, 3.645324e-14, 3.64262e-14, 3.66096e-14, 
    3.654319e-14, 3.672193e-14, 3.667367e-14, 3.675273e-14, 3.671345e-14, 
    3.670767e-14, 3.66572e-14, 3.662575e-14, 3.654624e-14, 3.648149e-14, 
    3.643012e-14, 3.644207e-14, 3.649849e-14, 3.660057e-14, 3.669705e-14, 
    3.667592e-14, 3.674673e-14, 3.655922e-14, 3.663788e-14, 3.660748e-14, 
    3.668674e-14, 3.6513e-14, 3.666087e-14, 3.647514e-14, 3.649145e-14, 
    3.654188e-14, 3.664319e-14, 3.666564e-14, 3.668954e-14, 3.66748e-14, 
    3.660317e-14, 3.659144e-14, 3.654066e-14, 3.652662e-14, 3.64879e-14, 
    3.645582e-14, 3.648512e-14, 3.651588e-14, 3.660321e-14, 3.668181e-14, 
    3.676742e-14, 3.678837e-14, 3.688816e-14, 3.680689e-14, 3.694091e-14, 
    3.682692e-14, 3.702417e-14, 3.666948e-14, 3.682363e-14, 3.654418e-14, 
    3.657434e-14, 3.662884e-14, 3.675374e-14, 3.668637e-14, 3.676517e-14, 
    3.659098e-14, 3.650041e-14, 3.647701e-14, 3.643324e-14, 3.647801e-14, 
    3.647437e-14, 3.651718e-14, 3.650342e-14, 3.660611e-14, 3.655097e-14, 
    3.670752e-14, 3.676455e-14, 3.692544e-14, 3.702386e-14, 3.712397e-14, 
    3.71681e-14, 3.718153e-14, 3.718715e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.200402e-14, 1.203457e-14, 1.202864e-14, 1.205326e-14, 1.203961e-14, 
    1.205572e-14, 1.201022e-14, 1.203578e-14, 1.201947e-14, 1.200677e-14, 
    1.210096e-14, 1.205436e-14, 1.214933e-14, 1.211966e-14, 1.219413e-14, 
    1.214471e-14, 1.220408e-14, 1.219272e-14, 1.222695e-14, 1.221714e-14, 
    1.226085e-14, 1.223147e-14, 1.22835e-14, 1.225384e-14, 1.225848e-14, 
    1.22305e-14, 1.206375e-14, 1.209516e-14, 1.206189e-14, 1.206637e-14, 
    1.206436e-14, 1.203988e-14, 1.202753e-14, 1.200169e-14, 1.200638e-14, 
    1.202537e-14, 1.206838e-14, 1.20538e-14, 1.209057e-14, 1.208974e-14, 
    1.21306e-14, 1.211218e-14, 1.218078e-14, 1.216131e-14, 1.221755e-14, 
    1.220342e-14, 1.221689e-14, 1.221281e-14, 1.221694e-14, 1.219621e-14, 
    1.220509e-14, 1.218684e-14, 1.211563e-14, 1.213658e-14, 1.207405e-14, 
    1.203637e-14, 1.201134e-14, 1.199355e-14, 1.199607e-14, 1.200086e-14, 
    1.202548e-14, 1.204862e-14, 1.206624e-14, 1.207802e-14, 1.208962e-14, 
    1.212467e-14, 1.214323e-14, 1.218471e-14, 1.217724e-14, 1.218991e-14, 
    1.220201e-14, 1.222231e-14, 1.221897e-14, 1.222791e-14, 1.218958e-14, 
    1.221506e-14, 1.217298e-14, 1.21845e-14, 1.209273e-14, 1.205774e-14, 
    1.204282e-14, 1.202978e-14, 1.1998e-14, 1.201995e-14, 1.20113e-14, 
    1.203188e-14, 1.204494e-14, 1.203848e-14, 1.207834e-14, 1.206285e-14, 
    1.214433e-14, 1.210926e-14, 1.22006e-14, 1.217878e-14, 1.220583e-14, 
    1.219203e-14, 1.221567e-14, 1.21944e-14, 1.223124e-14, 1.223925e-14, 
    1.223378e-14, 1.225481e-14, 1.219321e-14, 1.221688e-14, 1.20383e-14, 
    1.203935e-14, 1.204427e-14, 1.202267e-14, 1.202135e-14, 1.200155e-14, 
    1.201917e-14, 1.202667e-14, 1.20457e-14, 1.205695e-14, 1.206764e-14, 
    1.209112e-14, 1.211732e-14, 1.215392e-14, 1.218019e-14, 1.219778e-14, 
    1.2187e-14, 1.219652e-14, 1.218588e-14, 1.218089e-14, 1.223625e-14, 
    1.220517e-14, 1.225179e-14, 1.224921e-14, 1.222812e-14, 1.22495e-14, 
    1.204009e-14, 1.203403e-14, 1.201296e-14, 1.202945e-14, 1.19994e-14, 
    1.201622e-14, 1.202588e-14, 1.206317e-14, 1.207136e-14, 1.207894e-14, 
    1.209392e-14, 1.211313e-14, 1.214678e-14, 1.217604e-14, 1.220272e-14, 
    1.220077e-14, 1.220145e-14, 1.22074e-14, 1.219265e-14, 1.220983e-14, 
    1.22127e-14, 1.220517e-14, 1.224887e-14, 1.223639e-14, 1.224916e-14, 
    1.224104e-14, 1.2036e-14, 1.204621e-14, 1.204069e-14, 1.205106e-14, 
    1.204375e-14, 1.207621e-14, 1.208593e-14, 1.213138e-14, 1.211275e-14, 
    1.214241e-14, 1.211576e-14, 1.212049e-14, 1.214336e-14, 1.211721e-14, 
    1.217442e-14, 1.213563e-14, 1.220764e-14, 1.216894e-14, 1.221006e-14, 
    1.22026e-14, 1.221495e-14, 1.2226e-14, 1.22399e-14, 1.226552e-14, 
    1.225959e-14, 1.2281e-14, 1.206141e-14, 1.207463e-14, 1.207347e-14, 
    1.20873e-14, 1.209752e-14, 1.211967e-14, 1.215515e-14, 1.214182e-14, 
    1.21663e-14, 1.217121e-14, 1.213402e-14, 1.215685e-14, 1.208348e-14, 
    1.209534e-14, 1.208828e-14, 1.206245e-14, 1.214488e-14, 1.210261e-14, 
    1.218062e-14, 1.215776e-14, 1.222442e-14, 1.219129e-14, 1.225632e-14, 
    1.228405e-14, 1.231016e-14, 1.234059e-14, 1.208185e-14, 1.207287e-14, 
    1.208895e-14, 1.211117e-14, 1.213178e-14, 1.215916e-14, 1.216196e-14, 
    1.216708e-14, 1.218035e-14, 1.21915e-14, 1.216869e-14, 1.21943e-14, 
    1.209807e-14, 1.214855e-14, 1.206947e-14, 1.20933e-14, 1.210986e-14, 
    1.21026e-14, 1.21403e-14, 1.214917e-14, 1.218519e-14, 1.216658e-14, 
    1.227721e-14, 1.222832e-14, 1.236376e-14, 1.232598e-14, 1.206973e-14, 
    1.208182e-14, 1.212384e-14, 1.210386e-14, 1.216099e-14, 1.217503e-14, 
    1.218644e-14, 1.220101e-14, 1.220259e-14, 1.221122e-14, 1.219708e-14, 
    1.221066e-14, 1.215921e-14, 1.218222e-14, 1.211905e-14, 1.213444e-14, 
    1.212736e-14, 1.211959e-14, 1.214356e-14, 1.216905e-14, 1.216961e-14, 
    1.217777e-14, 1.220076e-14, 1.216122e-14, 1.228349e-14, 1.220803e-14, 
    1.209499e-14, 1.211824e-14, 1.212157e-14, 1.211257e-14, 1.217362e-14, 
    1.215151e-14, 1.221101e-14, 1.219495e-14, 1.222126e-14, 1.220819e-14, 
    1.220626e-14, 1.218946e-14, 1.217899e-14, 1.215253e-14, 1.213097e-14, 
    1.211387e-14, 1.211785e-14, 1.213663e-14, 1.217061e-14, 1.220273e-14, 
    1.219569e-14, 1.221927e-14, 1.215685e-14, 1.218303e-14, 1.217291e-14, 
    1.21993e-14, 1.214146e-14, 1.219069e-14, 1.212886e-14, 1.213429e-14, 
    1.215107e-14, 1.21848e-14, 1.219227e-14, 1.220023e-14, 1.219532e-14, 
    1.217148e-14, 1.216757e-14, 1.215067e-14, 1.214599e-14, 1.213311e-14, 
    1.212243e-14, 1.213218e-14, 1.214242e-14, 1.217149e-14, 1.219766e-14, 
    1.222615e-14, 1.223313e-14, 1.226635e-14, 1.223929e-14, 1.22839e-14, 
    1.224596e-14, 1.231162e-14, 1.219355e-14, 1.224486e-14, 1.215184e-14, 
    1.216188e-14, 1.218002e-14, 1.22216e-14, 1.219917e-14, 1.22254e-14, 
    1.216742e-14, 1.213727e-14, 1.212948e-14, 1.211491e-14, 1.212981e-14, 
    1.21286e-14, 1.214285e-14, 1.213828e-14, 1.217246e-14, 1.21541e-14, 
    1.220621e-14, 1.22252e-14, 1.227875e-14, 1.231152e-14, 1.234484e-14, 
    1.235954e-14, 1.236401e-14, 1.236587e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -1.003379e-10, -1.006127e-10, -1.005593e-10, -1.00781e-10, -1.00658e-10, 
    -1.008032e-10, -1.003936e-10, -1.006236e-10, -1.004768e-10, 
    -1.003626e-10, -1.012109e-10, -1.007909e-10, -1.016472e-10, 
    -1.013794e-10, -1.020521e-10, -1.016056e-10, -1.021421e-10, 
    -1.020393e-10, -1.023489e-10, -1.022602e-10, -1.026561e-10, 
    -1.023898e-10, -1.028613e-10, -1.025925e-10, -1.026346e-10, -1.02381e-10, 
    -1.008754e-10, -1.011586e-10, -1.008587e-10, -1.00899e-10, -1.008809e-10, 
    -1.006606e-10, -1.005495e-10, -1.003169e-10, -1.003591e-10, -1.0053e-10, 
    -1.009172e-10, -1.007858e-10, -1.01117e-10, -1.011096e-10, -1.014782e-10, 
    -1.01312e-10, -1.019314e-10, -1.017554e-10, -1.022639e-10, -1.02136e-10, 
    -1.022579e-10, -1.02221e-10, -1.022584e-10, -1.020708e-10, -1.021512e-10, 
    -1.019862e-10, -1.013431e-10, -1.015321e-10, -1.009682e-10, -1.00629e-10, 
    -1.004037e-10, -1.002438e-10, -1.002664e-10, -1.003095e-10, -1.00531e-10, 
    -1.007392e-10, -1.008978e-10, -1.010039e-10, -1.011085e-10, 
    -1.014247e-10, -1.015922e-10, -1.019669e-10, -1.018994e-10, 
    -1.020139e-10, -1.021233e-10, -1.02307e-10, -1.022768e-10, -1.023577e-10, 
    -1.020109e-10, -1.022414e-10, -1.018609e-10, -1.019649e-10, 
    -1.011368e-10, -1.008213e-10, -1.00687e-10, -1.005696e-10, -1.002838e-10, 
    -1.004811e-10, -1.004033e-10, -1.005885e-10, -1.007061e-10, 
    -1.006479e-10, -1.010068e-10, -1.008673e-10, -1.016021e-10, 
    -1.012857e-10, -1.021105e-10, -1.019132e-10, -1.021578e-10, -1.02033e-10, 
    -1.022469e-10, -1.020544e-10, -1.023878e-10, -1.024603e-10, 
    -1.024108e-10, -1.026013e-10, -1.020438e-10, -1.022579e-10, 
    -1.006463e-10, -1.006558e-10, -1.007e-10, -1.005057e-10, -1.004938e-10, 
    -1.003157e-10, -1.004742e-10, -1.005416e-10, -1.007129e-10, 
    -1.008142e-10, -1.009104e-10, -1.011221e-10, -1.013584e-10, 
    -1.016887e-10, -1.01926e-10, -1.02085e-10, -1.019876e-10, -1.020736e-10, 
    -1.019774e-10, -1.019323e-10, -1.024331e-10, -1.021519e-10, 
    -1.025739e-10, -1.025505e-10, -1.023596e-10, -1.025532e-10, 
    -1.006624e-10, -1.006078e-10, -1.004183e-10, -1.005666e-10, 
    -1.002963e-10, -1.004476e-10, -1.005346e-10, -1.008702e-10, 
    -1.009439e-10, -1.010123e-10, -1.011473e-10, -1.013205e-10, 
    -1.016243e-10, -1.018885e-10, -1.021297e-10, -1.02112e-10, -1.021182e-10, 
    -1.021721e-10, -1.020387e-10, -1.02194e-10, -1.022201e-10, -1.021519e-10, 
    -1.025474e-10, -1.024344e-10, -1.0255e-10, -1.024765e-10, -1.006256e-10, 
    -1.007174e-10, -1.006678e-10, -1.007611e-10, -1.006954e-10, 
    -1.009877e-10, -1.010753e-10, -1.014853e-10, -1.013171e-10, 
    -1.015848e-10, -1.013443e-10, -1.013869e-10, -1.015934e-10, 
    -1.013573e-10, -1.018739e-10, -1.015236e-10, -1.021742e-10, 
    -1.018245e-10, -1.021961e-10, -1.021286e-10, -1.022403e-10, 
    -1.023404e-10, -1.024662e-10, -1.026983e-10, -1.026445e-10, 
    -1.028386e-10, -1.008544e-10, -1.009734e-10, -1.00963e-10, -1.010876e-10, 
    -1.011798e-10, -1.013795e-10, -1.016998e-10, -1.015794e-10, 
    -1.018005e-10, -1.018448e-10, -1.01509e-10, -1.017152e-10, -1.010532e-10, 
    -1.011601e-10, -1.010965e-10, -1.008637e-10, -1.016071e-10, 
    -1.012257e-10, -1.019299e-10, -1.017234e-10, -1.023261e-10, 
    -1.020264e-10, -1.02615e-10, -1.028664e-10, -1.031031e-10, -1.033795e-10, 
    -1.010385e-10, -1.009576e-10, -1.011025e-10, -1.013028e-10, 
    -1.014888e-10, -1.01736e-10, -1.017613e-10, -1.018076e-10, -1.019275e-10, 
    -1.020283e-10, -1.018222e-10, -1.020535e-10, -1.011849e-10, 
    -1.016402e-10, -1.009269e-10, -1.011417e-10, -1.01291e-10, -1.012256e-10, 
    -1.015656e-10, -1.016458e-10, -1.019713e-10, -1.01803e-10, -1.028043e-10, 
    -1.023614e-10, -1.0359e-10, -1.032468e-10, -1.009293e-10, -1.010382e-10, 
    -1.014172e-10, -1.012369e-10, -1.017525e-10, -1.018794e-10, 
    -1.019825e-10, -1.021143e-10, -1.021285e-10, -1.022066e-10, 
    -1.020787e-10, -1.022016e-10, -1.017365e-10, -1.019444e-10, 
    -1.013739e-10, -1.015128e-10, -1.014489e-10, -1.013788e-10, 
    -1.015951e-10, -1.018254e-10, -1.018304e-10, -1.019042e-10, 
    -1.021122e-10, -1.017546e-10, -1.028614e-10, -1.021779e-10, -1.01157e-10, 
    -1.013667e-10, -1.013967e-10, -1.013154e-10, -1.018666e-10, 
    -1.016669e-10, -1.022047e-10, -1.020594e-10, -1.022975e-10, 
    -1.021792e-10, -1.021618e-10, -1.020098e-10, -1.019152e-10, 
    -1.016761e-10, -1.014815e-10, -1.013272e-10, -1.013631e-10, 
    -1.015326e-10, -1.018395e-10, -1.021298e-10, -1.020662e-10, 
    -1.022794e-10, -1.017151e-10, -1.019517e-10, -1.018603e-10, 
    -1.020988e-10, -1.015762e-10, -1.020211e-10, -1.014624e-10, 
    -1.015114e-10, -1.01663e-10, -1.019678e-10, -1.020352e-10, -1.021072e-10, 
    -1.020628e-10, -1.018473e-10, -1.01812e-10, -1.016593e-10, -1.016171e-10, 
    -1.015008e-10, -1.014044e-10, -1.014924e-10, -1.015849e-10, 
    -1.018474e-10, -1.020839e-10, -1.023418e-10, -1.024049e-10, 
    -1.027059e-10, -1.024608e-10, -1.028652e-10, -1.025213e-10, 
    -1.031166e-10, -1.020469e-10, -1.025113e-10, -1.016699e-10, 
    -1.017606e-10, -1.019245e-10, -1.023006e-10, -1.020976e-10, -1.02335e-10, 
    -1.018106e-10, -1.015384e-10, -1.01468e-10, -1.013366e-10, -1.01471e-10, 
    -1.014601e-10, -1.015887e-10, -1.015474e-10, -1.018561e-10, 
    -1.016903e-10, -1.021613e-10, -1.023331e-10, -1.028183e-10, 
    -1.031155e-10, -1.034181e-10, -1.035516e-10, -1.035923e-10, -1.036093e-10 ;

 SMINN_TO_SOIL1N_S3 =
  -2.418215e-12, -2.424838e-12, -2.423551e-12, -2.428892e-12, -2.42593e-12, 
    -2.429426e-12, -2.419559e-12, -2.425101e-12, -2.421563e-12, 
    -2.418812e-12, -2.439251e-12, -2.42913e-12, -2.449764e-12, -2.443312e-12, 
    -2.459518e-12, -2.44876e-12, -2.461687e-12, -2.459209e-12, -2.46667e-12, 
    -2.464533e-12, -2.474071e-12, -2.467656e-12, -2.479015e-12, -2.47254e-12, 
    -2.473552e-12, -2.467444e-12, -2.431168e-12, -2.437991e-12, 
    -2.430763e-12, -2.431736e-12, -2.4313e-12, -2.42599e-12, -2.423314e-12, 
    -2.41771e-12, -2.418727e-12, -2.422844e-12, -2.432174e-12, -2.429008e-12, 
    -2.436989e-12, -2.436809e-12, -2.44569e-12, -2.441686e-12, -2.45661e-12, 
    -2.452369e-12, -2.464622e-12, -2.461541e-12, -2.464477e-12, 
    -2.463587e-12, -2.464488e-12, -2.45997e-12, -2.461906e-12, -2.45793e-12, 
    -2.442436e-12, -2.44699e-12, -2.433404e-12, -2.42523e-12, -2.419802e-12, 
    -2.415948e-12, -2.416493e-12, -2.417531e-12, -2.422868e-12, 
    -2.427885e-12, -2.431707e-12, -2.434264e-12, -2.436783e-12, 
    -2.444403e-12, -2.448437e-12, -2.457467e-12, -2.455838e-12, 
    -2.458597e-12, -2.461234e-12, -2.46566e-12, -2.464932e-12, -2.466881e-12, 
    -2.458525e-12, -2.464078e-12, -2.45491e-12, -2.457418e-12, -2.437464e-12, 
    -2.429862e-12, -2.426627e-12, -2.423799e-12, -2.416912e-12, 
    -2.421667e-12, -2.419793e-12, -2.424254e-12, -2.427087e-12, 
    -2.425686e-12, -2.434334e-12, -2.430972e-12, -2.448676e-12, 
    -2.441052e-12, -2.460927e-12, -2.456173e-12, -2.462066e-12, 
    -2.459059e-12, -2.464211e-12, -2.459575e-12, -2.467607e-12, 
    -2.469355e-12, -2.46816e-12, -2.47275e-12, -2.459317e-12, -2.464477e-12, 
    -2.425646e-12, -2.425875e-12, -2.42694e-12, -2.422258e-12, -2.421972e-12, 
    -2.417682e-12, -2.421499e-12, -2.423125e-12, -2.427252e-12, 
    -2.429692e-12, -2.432011e-12, -2.43711e-12, -2.442804e-12, -2.450763e-12, 
    -2.456481e-12, -2.460312e-12, -2.457963e-12, -2.460037e-12, 
    -2.457718e-12, -2.456632e-12, -2.4687e-12, -2.461924e-12, -2.47209e-12, 
    -2.471528e-12, -2.466927e-12, -2.471591e-12, -2.426035e-12, -2.42472e-12, 
    -2.420153e-12, -2.423727e-12, -2.417214e-12, -2.42086e-12, -2.422955e-12, 
    -2.431041e-12, -2.432818e-12, -2.434465e-12, -2.437718e-12, 
    -2.441891e-12, -2.44921e-12, -2.455577e-12, -2.461388e-12, -2.460962e-12, 
    -2.461112e-12, -2.46241e-12, -2.459195e-12, -2.462938e-12, -2.463565e-12, 
    -2.461923e-12, -2.471453e-12, -2.468731e-12, -2.471516e-12, 
    -2.469744e-12, -2.425148e-12, -2.427361e-12, -2.426165e-12, 
    -2.428413e-12, -2.426829e-12, -2.433872e-12, -2.435983e-12, 
    -2.445861e-12, -2.441809e-12, -2.448259e-12, -2.442464e-12, 
    -2.443491e-12, -2.448468e-12, -2.442778e-12, -2.455225e-12, 
    -2.446786e-12, -2.46246e-12, -2.454034e-12, -2.462988e-12, -2.461363e-12, 
    -2.464054e-12, -2.466464e-12, -2.469496e-12, -2.475088e-12, 
    -2.473793e-12, -2.478469e-12, -2.43066e-12, -2.433529e-12, -2.433277e-12, 
    -2.43628e-12, -2.438501e-12, -2.443314e-12, -2.45103e-12, -2.448129e-12, 
    -2.453456e-12, -2.454525e-12, -2.446432e-12, -2.451401e-12, -2.43545e-12, 
    -2.438027e-12, -2.436493e-12, -2.430886e-12, -2.448797e-12, 
    -2.439606e-12, -2.456575e-12, -2.451598e-12, -2.46612e-12, -2.458899e-12, 
    -2.47308e-12, -2.479138e-12, -2.484842e-12, -2.491502e-12, -2.435096e-12, 
    -2.433146e-12, -2.436637e-12, -2.441466e-12, -2.445947e-12, 
    -2.451902e-12, -2.452512e-12, -2.453627e-12, -2.456516e-12, 
    -2.458945e-12, -2.453979e-12, -2.459553e-12, -2.438623e-12, 
    -2.449594e-12, -2.432409e-12, -2.437584e-12, -2.441182e-12, 
    -2.439604e-12, -2.447798e-12, -2.449728e-12, -2.457571e-12, 
    -2.453517e-12, -2.477643e-12, -2.466972e-12, -2.496574e-12, 
    -2.488304e-12, -2.432465e-12, -2.435089e-12, -2.444221e-12, 
    -2.439877e-12, -2.4523e-12, -2.455356e-12, -2.457841e-12, -2.461017e-12, 
    -2.46136e-12, -2.463241e-12, -2.460158e-12, -2.46312e-12, -2.451915e-12, 
    -2.456923e-12, -2.443178e-12, -2.446524e-12, -2.444985e-12, 
    -2.443296e-12, -2.448507e-12, -2.454056e-12, -2.454176e-12, 
    -2.455955e-12, -2.460965e-12, -2.45235e-12, -2.479017e-12, -2.46255e-12, 
    -2.437951e-12, -2.443003e-12, -2.443726e-12, -2.441769e-12, -2.45505e-12, 
    -2.450239e-12, -2.463195e-12, -2.459695e-12, -2.465431e-12, -2.46258e-12, 
    -2.462161e-12, -2.4585e-12, -2.45622e-12, -2.450459e-12, -2.445771e-12, 
    -2.442053e-12, -2.442918e-12, -2.447001e-12, -2.454396e-12, 
    -2.461391e-12, -2.459858e-12, -2.464995e-12, -2.451399e-12, -2.4571e-12, 
    -2.454897e-12, -2.460643e-12, -2.448052e-12, -2.458771e-12, -2.44531e-12, 
    -2.446491e-12, -2.450143e-12, -2.457486e-12, -2.459112e-12, 
    -2.460846e-12, -2.459777e-12, -2.454584e-12, -2.453734e-12, 
    -2.450054e-12, -2.449038e-12, -2.446234e-12, -2.443912e-12, 
    -2.446034e-12, -2.448261e-12, -2.454587e-12, -2.460286e-12, 
    -2.466498e-12, -2.468018e-12, -2.475271e-12, -2.469366e-12, 
    -2.479109e-12, -2.470824e-12, -2.485166e-12, -2.459394e-12, 
    -2.470582e-12, -2.450309e-12, -2.452495e-12, -2.456445e-12, 
    -2.465506e-12, -2.460616e-12, -2.466335e-12, -2.453701e-12, 
    -2.447142e-12, -2.445446e-12, -2.442279e-12, -2.445518e-12, 
    -2.445255e-12, -2.448354e-12, -2.447358e-12, -2.454797e-12, 
    -2.450801e-12, -2.46215e-12, -2.46629e-12, -2.477979e-12, -2.485141e-12, 
    -2.492431e-12, -2.495649e-12, -2.496628e-12, -2.497037e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.899552e-15, 3.909478e-15, 3.907551e-15, 3.915549e-15, 3.911114e-15, 
    3.916349e-15, 3.901567e-15, 3.909871e-15, 3.904572e-15, 3.900448e-15, 
    3.931045e-15, 3.915906e-15, 3.946757e-15, 3.93712e-15, 3.961311e-15, 
    3.945256e-15, 3.964545e-15, 3.960852e-15, 3.971972e-15, 3.968788e-15, 
    3.982987e-15, 3.973441e-15, 3.990343e-15, 3.98071e-15, 3.982217e-15, 
    3.973125e-15, 3.918958e-15, 3.92916e-15, 3.918352e-15, 3.919808e-15, 
    3.919156e-15, 3.911205e-15, 3.907193e-15, 3.898795e-15, 3.900321e-15, 
    3.90649e-15, 3.920463e-15, 3.915724e-15, 3.927668e-15, 3.927399e-15, 
    3.940674e-15, 3.934691e-15, 3.956976e-15, 3.950649e-15, 3.968921e-15, 
    3.964329e-15, 3.968705e-15, 3.967379e-15, 3.968722e-15, 3.961987e-15, 
    3.964873e-15, 3.958945e-15, 3.935811e-15, 3.942616e-15, 3.922304e-15, 
    3.910062e-15, 3.901931e-15, 3.896153e-15, 3.89697e-15, 3.898527e-15, 
    3.906526e-15, 3.914043e-15, 3.919766e-15, 3.923592e-15, 3.92736e-15, 
    3.938747e-15, 3.944776e-15, 3.958253e-15, 3.955825e-15, 3.95994e-15, 
    3.963872e-15, 3.970467e-15, 3.969382e-15, 3.972286e-15, 3.959833e-15, 
    3.96811e-15, 3.954442e-15, 3.958182e-15, 3.928372e-15, 3.917003e-15, 
    3.912156e-15, 3.907921e-15, 3.897598e-15, 3.904727e-15, 3.901917e-15, 
    3.908603e-15, 3.912848e-15, 3.910749e-15, 3.923696e-15, 3.918665e-15, 
    3.945133e-15, 3.933743e-15, 3.963414e-15, 3.956324e-15, 3.965113e-15, 
    3.96063e-15, 3.968309e-15, 3.961398e-15, 3.973367e-15, 3.97597e-15, 
    3.974191e-15, 3.981025e-15, 3.961014e-15, 3.968704e-15, 3.91069e-15, 
    3.911032e-15, 3.912628e-15, 3.905612e-15, 3.905184e-15, 3.898753e-15, 
    3.904476e-15, 3.906911e-15, 3.913095e-15, 3.916748e-15, 3.92022e-15, 
    3.927849e-15, 3.93636e-15, 3.94825e-15, 3.956784e-15, 3.962498e-15, 
    3.958995e-15, 3.962088e-15, 3.95863e-15, 3.95701e-15, 3.974993e-15, 
    3.964899e-15, 3.980043e-15, 3.979206e-15, 3.972355e-15, 3.9793e-15, 
    3.911272e-15, 3.909303e-15, 3.902457e-15, 3.907815e-15, 3.898052e-15, 
    3.903517e-15, 3.906657e-15, 3.918767e-15, 3.921429e-15, 3.923892e-15, 
    3.928758e-15, 3.934997e-15, 3.945931e-15, 3.955434e-15, 3.964101e-15, 
    3.963467e-15, 3.96369e-15, 3.965624e-15, 3.960832e-15, 3.966411e-15, 
    3.967346e-15, 3.964899e-15, 3.979094e-15, 3.975041e-15, 3.979188e-15, 
    3.97655e-15, 3.909943e-15, 3.913258e-15, 3.911467e-15, 3.914834e-15, 
    3.912461e-15, 3.923003e-15, 3.926162e-15, 3.940928e-15, 3.934874e-15, 
    3.94451e-15, 3.935854e-15, 3.937388e-15, 3.944819e-15, 3.936323e-15, 
    3.954908e-15, 3.942308e-15, 3.965699e-15, 3.953129e-15, 3.966486e-15, 
    3.964064e-15, 3.968075e-15, 3.971665e-15, 3.97618e-15, 3.984502e-15, 
    3.982576e-15, 3.989532e-15, 3.918198e-15, 3.922491e-15, 3.922115e-15, 
    3.926608e-15, 3.929929e-15, 3.937124e-15, 3.948649e-15, 3.944318e-15, 
    3.952271e-15, 3.953865e-15, 3.941784e-15, 3.949202e-15, 3.925365e-15, 
    3.929219e-15, 3.926926e-15, 3.918535e-15, 3.945313e-15, 3.93158e-15, 
    3.956924e-15, 3.949498e-15, 3.971153e-15, 3.960388e-15, 3.981515e-15, 
    3.990524e-15, 3.999004e-15, 4.008889e-15, 3.924836e-15, 3.921919e-15, 
    3.927143e-15, 3.93436e-15, 3.941058e-15, 3.949951e-15, 3.950861e-15, 
    3.952525e-15, 3.956836e-15, 3.960459e-15, 3.953049e-15, 3.961366e-15, 
    3.930107e-15, 3.946505e-15, 3.920814e-15, 3.928555e-15, 3.933936e-15, 
    3.931578e-15, 3.943824e-15, 3.946706e-15, 3.958409e-15, 3.952362e-15, 
    3.9883e-15, 3.972419e-15, 4.016416e-15, 4.004144e-15, 3.920899e-15, 
    3.924827e-15, 3.938478e-15, 3.931986e-15, 3.950545e-15, 3.955106e-15, 
    3.958814e-15, 3.963547e-15, 3.96406e-15, 3.966863e-15, 3.962269e-15, 
    3.966683e-15, 3.94997e-15, 3.957443e-15, 3.936921e-15, 3.94192e-15, 
    3.939621e-15, 3.937099e-15, 3.944883e-15, 3.953165e-15, 3.953345e-15, 
    3.955999e-15, 3.963464e-15, 3.95062e-15, 3.99034e-15, 3.965827e-15, 
    3.929107e-15, 3.936658e-15, 3.937741e-15, 3.934816e-15, 3.954649e-15, 
    3.947467e-15, 3.966795e-15, 3.961577e-15, 3.970126e-15, 3.965879e-15, 
    3.965254e-15, 3.959796e-15, 3.956394e-15, 3.947796e-15, 3.940795e-15, 
    3.935241e-15, 3.936533e-15, 3.942633e-15, 3.953672e-15, 3.964104e-15, 
    3.96182e-15, 3.969477e-15, 3.9492e-15, 3.957707e-15, 3.954419e-15, 
    3.96299e-15, 3.944202e-15, 3.960193e-15, 3.940108e-15, 3.941872e-15, 
    3.947325e-15, 3.958281e-15, 3.960709e-15, 3.963293e-15, 3.961699e-15, 
    3.953953e-15, 3.952685e-15, 3.947193e-15, 3.945675e-15, 3.941488e-15, 
    3.938019e-15, 3.941188e-15, 3.944514e-15, 3.953958e-15, 3.962457e-15, 
    3.971715e-15, 3.97398e-15, 3.984772e-15, 3.975983e-15, 3.990475e-15, 
    3.978148e-15, 3.999479e-15, 3.961124e-15, 3.977793e-15, 3.947574e-15, 
    3.950836e-15, 3.956728e-15, 3.970235e-15, 3.96295e-15, 3.971471e-15, 
    3.952635e-15, 3.942841e-15, 3.94031e-15, 3.935578e-15, 3.940418e-15, 
    3.940025e-15, 3.944654e-15, 3.943167e-15, 3.954271e-15, 3.948309e-15, 
    3.965237e-15, 3.971405e-15, 3.988802e-15, 3.999446e-15, 4.010272e-15, 
    4.015044e-15, 4.016497e-15, 4.017104e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -1.050255e-08, -1.053129e-08, -1.052571e-08, -1.054889e-08, -1.053603e-08, 
    -1.055121e-08, -1.050838e-08, -1.053243e-08, -1.051708e-08, 
    -1.050514e-08, -1.059384e-08, -1.054992e-08, -1.063947e-08, 
    -1.061147e-08, -1.06818e-08, -1.063511e-08, -1.069122e-08, -1.068046e-08, 
    -1.071284e-08, -1.070357e-08, -1.074496e-08, -1.071712e-08, 
    -1.076642e-08, -1.073832e-08, -1.074271e-08, -1.07162e-08, -1.055877e-08, 
    -1.058838e-08, -1.055701e-08, -1.056123e-08, -1.055934e-08, -1.05363e-08, 
    -1.052468e-08, -1.050036e-08, -1.050477e-08, -1.052264e-08, 
    -1.056313e-08, -1.054939e-08, -1.058403e-08, -1.058325e-08, 
    -1.062179e-08, -1.060441e-08, -1.066918e-08, -1.065078e-08, 
    -1.070395e-08, -1.069058e-08, -1.070333e-08, -1.069946e-08, 
    -1.070338e-08, -1.068376e-08, -1.069217e-08, -1.067491e-08, 
    -1.060767e-08, -1.062743e-08, -1.056847e-08, -1.053299e-08, 
    -1.050944e-08, -1.049271e-08, -1.049508e-08, -1.049958e-08, 
    -1.052274e-08, -1.054452e-08, -1.056111e-08, -1.05722e-08, -1.058313e-08, 
    -1.06162e-08, -1.063371e-08, -1.06729e-08, -1.066583e-08, -1.067781e-08, 
    -1.068925e-08, -1.070846e-08, -1.07053e-08, -1.071376e-08, -1.06775e-08, 
    -1.07016e-08, -1.066181e-08, -1.067269e-08, -1.058609e-08, -1.05531e-08, 
    -1.053906e-08, -1.052678e-08, -1.049689e-08, -1.051753e-08, -1.05094e-08, 
    -1.052876e-08, -1.054105e-08, -1.053497e-08, -1.05725e-08, -1.055791e-08, 
    -1.063475e-08, -1.060166e-08, -1.068792e-08, -1.066728e-08, 
    -1.069286e-08, -1.067981e-08, -1.070217e-08, -1.068205e-08, 
    -1.071691e-08, -1.07245e-08, -1.071931e-08, -1.073923e-08, -1.068093e-08, 
    -1.070332e-08, -1.05348e-08, -1.053579e-08, -1.054041e-08, -1.05201e-08, 
    -1.051885e-08, -1.050024e-08, -1.05168e-08, -1.052386e-08, -1.054177e-08, 
    -1.055236e-08, -1.056242e-08, -1.058455e-08, -1.060926e-08, 
    -1.064381e-08, -1.066862e-08, -1.068525e-08, -1.067506e-08, 
    -1.068406e-08, -1.067399e-08, -1.066928e-08, -1.072165e-08, 
    -1.069225e-08, -1.073637e-08, -1.073393e-08, -1.071396e-08, -1.07342e-08, 
    -1.053649e-08, -1.053078e-08, -1.051096e-08, -1.052647e-08, 
    -1.049821e-08, -1.051403e-08, -1.052312e-08, -1.055822e-08, 
    -1.056593e-08, -1.057307e-08, -1.058719e-08, -1.06053e-08, -1.063707e-08, 
    -1.06647e-08, -1.068992e-08, -1.068807e-08, -1.068872e-08, -1.069435e-08, 
    -1.06804e-08, -1.069664e-08, -1.069937e-08, -1.069224e-08, -1.07336e-08, 
    -1.072179e-08, -1.073387e-08, -1.072618e-08, -1.053264e-08, 
    -1.054224e-08, -1.053705e-08, -1.054681e-08, -1.053994e-08, -1.05705e-08, 
    -1.057967e-08, -1.062253e-08, -1.060495e-08, -1.063294e-08, 
    -1.060779e-08, -1.061225e-08, -1.063385e-08, -1.060915e-08, 
    -1.066317e-08, -1.062654e-08, -1.069457e-08, -1.0658e-08, -1.069686e-08, 
    -1.068981e-08, -1.070149e-08, -1.071195e-08, -1.072511e-08, 
    -1.074937e-08, -1.074376e-08, -1.076405e-08, -1.055656e-08, 
    -1.056901e-08, -1.056792e-08, -1.058095e-08, -1.059059e-08, 
    -1.061148e-08, -1.064497e-08, -1.063238e-08, -1.065549e-08, 
    -1.066013e-08, -1.062501e-08, -1.064657e-08, -1.057735e-08, 
    -1.058853e-08, -1.058188e-08, -1.055754e-08, -1.063527e-08, 
    -1.059539e-08, -1.066903e-08, -1.064743e-08, -1.071046e-08, 
    -1.067912e-08, -1.074066e-08, -1.076695e-08, -1.079171e-08, 
    -1.082061e-08, -1.057581e-08, -1.056735e-08, -1.05825e-08, -1.060346e-08, 
    -1.062291e-08, -1.064875e-08, -1.06514e-08, -1.065624e-08, -1.066877e-08, 
    -1.067932e-08, -1.065776e-08, -1.068196e-08, -1.059112e-08, 
    -1.063874e-08, -1.056415e-08, -1.058661e-08, -1.060222e-08, 
    -1.059538e-08, -1.063094e-08, -1.063932e-08, -1.067335e-08, 
    -1.065576e-08, -1.076046e-08, -1.071415e-08, -1.084262e-08, 
    -1.080674e-08, -1.056439e-08, -1.057578e-08, -1.061541e-08, 
    -1.059656e-08, -1.065048e-08, -1.066374e-08, -1.067453e-08, 
    -1.068831e-08, -1.06898e-08, -1.069796e-08, -1.068458e-08, -1.069743e-08, 
    -1.06488e-08, -1.067054e-08, -1.061089e-08, -1.062541e-08, -1.061873e-08, 
    -1.06114e-08, -1.063402e-08, -1.06581e-08, -1.065862e-08, -1.066634e-08, 
    -1.068809e-08, -1.06507e-08, -1.076643e-08, -1.069496e-08, -1.05882e-08, 
    -1.061013e-08, -1.061327e-08, -1.060477e-08, -1.066241e-08, 
    -1.064153e-08, -1.069776e-08, -1.068257e-08, -1.070747e-08, 
    -1.069509e-08, -1.069327e-08, -1.067739e-08, -1.066749e-08, 
    -1.064249e-08, -1.062214e-08, -1.060601e-08, -1.060976e-08, 
    -1.062748e-08, -1.065958e-08, -1.068993e-08, -1.068328e-08, 
    -1.070557e-08, -1.064657e-08, -1.067131e-08, -1.066175e-08, 
    -1.068668e-08, -1.063204e-08, -1.067856e-08, -1.062014e-08, 
    -1.062527e-08, -1.064112e-08, -1.067299e-08, -1.068004e-08, 
    -1.068757e-08, -1.068293e-08, -1.066039e-08, -1.06567e-08, -1.064073e-08, 
    -1.063632e-08, -1.062415e-08, -1.061407e-08, -1.062328e-08, 
    -1.063295e-08, -1.06604e-08, -1.068514e-08, -1.07121e-08, -1.071869e-08, 
    -1.075017e-08, -1.072454e-08, -1.076683e-08, -1.073087e-08, 
    -1.079311e-08, -1.068126e-08, -1.072982e-08, -1.064184e-08, 
    -1.065132e-08, -1.066847e-08, -1.070779e-08, -1.068657e-08, 
    -1.071139e-08, -1.065656e-08, -1.062809e-08, -1.062073e-08, 
    -1.060699e-08, -1.062104e-08, -1.06199e-08, -1.063335e-08, -1.062903e-08, 
    -1.066131e-08, -1.064397e-08, -1.069323e-08, -1.071119e-08, 
    -1.076192e-08, -1.079301e-08, -1.082465e-08, -1.083861e-08, 
    -1.084286e-08, -1.084463e-08 ;

 SMINN_TO_SOIL3N_S1 =
  -1.246122e-10, -1.249534e-10, -1.248871e-10, -1.251622e-10, -1.250096e-10, 
    -1.251898e-10, -1.246814e-10, -1.249669e-10, -1.247847e-10, -1.24643e-10, 
    -1.256959e-10, -1.251745e-10, -1.262375e-10, -1.259051e-10, 
    -1.267401e-10, -1.261858e-10, -1.268518e-10, -1.267242e-10, 
    -1.271085e-10, -1.269984e-10, -1.274899e-10, -1.271594e-10, 
    -1.277446e-10, -1.27411e-10, -1.274631e-10, -1.271485e-10, -1.252795e-10, 
    -1.25631e-10, -1.252587e-10, -1.253088e-10, -1.252863e-10, -1.250128e-10, 
    -1.248749e-10, -1.245862e-10, -1.246386e-10, -1.248507e-10, 
    -1.253313e-10, -1.251682e-10, -1.255794e-10, -1.255701e-10, 
    -1.260277e-10, -1.258214e-10, -1.265903e-10, -1.263718e-10, -1.27003e-10, 
    -1.268443e-10, -1.269956e-10, -1.269497e-10, -1.269962e-10, 
    -1.267634e-10, -1.268631e-10, -1.266583e-10, -1.2586e-10, -1.260946e-10, 
    -1.253947e-10, -1.249736e-10, -1.246939e-10, -1.244954e-10, 
    -1.245235e-10, -1.24577e-10, -1.248519e-10, -1.251104e-10, -1.253073e-10, 
    -1.25439e-10, -1.255688e-10, -1.259613e-10, -1.261692e-10, -1.266344e-10, 
    -1.265505e-10, -1.266927e-10, -1.268285e-10, -1.270565e-10, -1.27019e-10, 
    -1.271194e-10, -1.26689e-10, -1.26975e-10, -1.265027e-10, -1.266319e-10, 
    -1.256039e-10, -1.252122e-10, -1.250456e-10, -1.248998e-10, 
    -1.245451e-10, -1.247901e-10, -1.246935e-10, -1.249233e-10, 
    -1.250693e-10, -1.249971e-10, -1.254426e-10, -1.252694e-10, 
    -1.261815e-10, -1.257887e-10, -1.268127e-10, -1.265677e-10, 
    -1.268714e-10, -1.267165e-10, -1.269819e-10, -1.26743e-10, -1.271568e-10, 
    -1.272469e-10, -1.271853e-10, -1.274218e-10, -1.267298e-10, 
    -1.269956e-10, -1.24995e-10, -1.250068e-10, -1.250617e-10, -1.248205e-10, 
    -1.248057e-10, -1.245847e-10, -1.247814e-10, -1.248651e-10, 
    -1.250777e-10, -1.252034e-10, -1.253229e-10, -1.255857e-10, -1.25879e-10, 
    -1.26289e-10, -1.265836e-10, -1.26781e-10, -1.2666e-10, -1.267668e-10, 
    -1.266474e-10, -1.265914e-10, -1.272131e-10, -1.26864e-10, -1.273878e-10, 
    -1.273588e-10, -1.271218e-10, -1.273621e-10, -1.250151e-10, 
    -1.249473e-10, -1.24712e-10, -1.248962e-10, -1.245607e-10, -1.247484e-10, 
    -1.248564e-10, -1.25273e-10, -1.253645e-10, -1.254494e-10, -1.256169e-10, 
    -1.258319e-10, -1.26209e-10, -1.26537e-10, -1.268364e-10, -1.268145e-10, 
    -1.268222e-10, -1.268891e-10, -1.267234e-10, -1.269163e-10, 
    -1.269486e-10, -1.26864e-10, -1.27355e-10, -1.272147e-10, -1.273582e-10, 
    -1.272669e-10, -1.249694e-10, -1.250834e-10, -1.250218e-10, 
    -1.251376e-10, -1.25056e-10, -1.254188e-10, -1.255276e-10, -1.260365e-10, 
    -1.258277e-10, -1.2616e-10, -1.258615e-10, -1.259144e-10, -1.261708e-10, 
    -1.258776e-10, -1.265189e-10, -1.260841e-10, -1.268917e-10, 
    -1.264575e-10, -1.269189e-10, -1.268351e-10, -1.269738e-10, 
    -1.270979e-10, -1.272541e-10, -1.275423e-10, -1.274755e-10, 
    -1.277165e-10, -1.252533e-10, -1.254012e-10, -1.253882e-10, 
    -1.255429e-10, -1.256573e-10, -1.259052e-10, -1.263028e-10, 
    -1.261533e-10, -1.264278e-10, -1.264828e-10, -1.260659e-10, 
    -1.263219e-10, -1.255001e-10, -1.256329e-10, -1.255538e-10, -1.25265e-10, 
    -1.261877e-10, -1.257142e-10, -1.265885e-10, -1.263321e-10, 
    -1.270802e-10, -1.267082e-10, -1.274388e-10, -1.277509e-10, 
    -1.280448e-10, -1.28388e-10, -1.254819e-10, -1.253814e-10, -1.255613e-10, 
    -1.2581e-10, -1.260409e-10, -1.263477e-10, -1.263791e-10, -1.264366e-10, 
    -1.265854e-10, -1.267105e-10, -1.264547e-10, -1.267419e-10, 
    -1.256636e-10, -1.262288e-10, -1.253434e-10, -1.256101e-10, 
    -1.257954e-10, -1.257141e-10, -1.261362e-10, -1.262357e-10, 
    -1.266398e-10, -1.264309e-10, -1.276739e-10, -1.271241e-10, 
    -1.286493e-10, -1.282232e-10, -1.253463e-10, -1.254815e-10, -1.25952e-10, 
    -1.257282e-10, -1.263682e-10, -1.265257e-10, -1.266537e-10, 
    -1.268173e-10, -1.26835e-10, -1.269319e-10, -1.267731e-10, -1.269257e-10, 
    -1.263483e-10, -1.266064e-10, -1.258983e-10, -1.260706e-10, 
    -1.259913e-10, -1.259043e-10, -1.261728e-10, -1.264587e-10, 
    -1.264649e-10, -1.265565e-10, -1.268147e-10, -1.263708e-10, 
    -1.277447e-10, -1.268963e-10, -1.25629e-10, -1.258893e-10, -1.259265e-10, 
    -1.258257e-10, -1.265099e-10, -1.26262e-10, -1.269296e-10, -1.267492e-10, 
    -1.270447e-10, -1.268979e-10, -1.268763e-10, -1.266876e-10, 
    -1.265702e-10, -1.262734e-10, -1.260318e-10, -1.258403e-10, 
    -1.258848e-10, -1.260952e-10, -1.264762e-10, -1.268366e-10, 
    -1.267576e-10, -1.270223e-10, -1.263218e-10, -1.266155e-10, -1.26502e-10, 
    -1.26798e-10, -1.261493e-10, -1.267016e-10, -1.260081e-10, -1.260689e-10, 
    -1.262571e-10, -1.266354e-10, -1.267192e-10, -1.268085e-10, 
    -1.267534e-10, -1.264859e-10, -1.264421e-10, -1.262525e-10, 
    -1.262001e-10, -1.260557e-10, -1.259361e-10, -1.260454e-10, 
    -1.261601e-10, -1.26486e-10, -1.267796e-10, -1.270997e-10, -1.27178e-10, 
    -1.275517e-10, -1.272475e-10, -1.277494e-10, -1.273226e-10, 
    -1.280615e-10, -1.267337e-10, -1.273101e-10, -1.262657e-10, 
    -1.263782e-10, -1.265818e-10, -1.270486e-10, -1.267966e-10, 
    -1.270913e-10, -1.264404e-10, -1.261025e-10, -1.260151e-10, 
    -1.258519e-10, -1.260188e-10, -1.260052e-10, -1.261649e-10, 
    -1.261136e-10, -1.264969e-10, -1.26291e-10, -1.268757e-10, -1.27089e-10, 
    -1.276912e-10, -1.280602e-10, -1.284358e-10, -1.286016e-10, 
    -1.286521e-10, -1.286732e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -1.033927e-11, -1.036759e-11, -1.036209e-11, -1.038492e-11, -1.037226e-11, 
    -1.038721e-11, -1.034501e-11, -1.036871e-11, -1.035358e-11, 
    -1.034182e-11, -1.042923e-11, -1.038594e-11, -1.047419e-11, 
    -1.044659e-11, -1.05159e-11, -1.046989e-11, -1.052518e-11, -1.051458e-11, 
    -1.054649e-11, -1.053735e-11, -1.057814e-11, -1.055071e-11, 
    -1.059929e-11, -1.05716e-11, -1.057593e-11, -1.05498e-11, -1.039466e-11, 
    -1.042384e-11, -1.039293e-11, -1.039709e-11, -1.039522e-11, 
    -1.037252e-11, -1.036107e-11, -1.03371e-11, -1.034145e-11, -1.035906e-11, 
    -1.039896e-11, -1.038542e-11, -1.041955e-11, -1.041878e-11, 
    -1.045677e-11, -1.043964e-11, -1.050347e-11, -1.048533e-11, 
    -1.053773e-11, -1.052456e-11, -1.053711e-11, -1.053331e-11, 
    -1.053716e-11, -1.051784e-11, -1.052612e-11, -1.050911e-11, 
    -1.044285e-11, -1.046233e-11, -1.040422e-11, -1.036926e-11, 
    -1.034605e-11, -1.032957e-11, -1.03319e-11, -1.033634e-11, -1.035916e-11, 
    -1.038062e-11, -1.039697e-11, -1.04079e-11, -1.041867e-11, -1.045126e-11, 
    -1.046852e-11, -1.050713e-11, -1.050017e-11, -1.051197e-11, 
    -1.052325e-11, -1.054217e-11, -1.053906e-11, -1.054739e-11, 
    -1.051166e-11, -1.053541e-11, -1.04962e-11, -1.050693e-11, -1.042159e-11, 
    -1.038908e-11, -1.037524e-11, -1.036314e-11, -1.033369e-11, 
    -1.035403e-11, -1.034601e-11, -1.036509e-11, -1.037721e-11, 
    -1.037121e-11, -1.04082e-11, -1.039382e-11, -1.046954e-11, -1.043693e-11, 
    -1.052193e-11, -1.05016e-11, -1.05268e-11, -1.051394e-11, -1.053598e-11, 
    -1.051615e-11, -1.05505e-11, -1.055797e-11, -1.055287e-11, -1.05725e-11, 
    -1.051505e-11, -1.053711e-11, -1.037105e-11, -1.037202e-11, 
    -1.037658e-11, -1.035655e-11, -1.035533e-11, -1.033698e-11, 
    -1.035331e-11, -1.036026e-11, -1.037791e-11, -1.038835e-11, 
    -1.039827e-11, -1.042007e-11, -1.044442e-11, -1.047846e-11, 
    -1.050292e-11, -1.05193e-11, -1.050926e-11, -1.051813e-11, -1.050821e-11, 
    -1.050356e-11, -1.055517e-11, -1.052619e-11, -1.056967e-11, 
    -1.056727e-11, -1.054759e-11, -1.056754e-11, -1.037271e-11, 
    -1.036708e-11, -1.034755e-11, -1.036284e-11, -1.033498e-11, 
    -1.035057e-11, -1.035954e-11, -1.039412e-11, -1.040172e-11, 
    -1.040876e-11, -1.042267e-11, -1.044052e-11, -1.047182e-11, 
    -1.049905e-11, -1.05239e-11, -1.052208e-11, -1.052272e-11, -1.052827e-11, 
    -1.051452e-11, -1.053053e-11, -1.053321e-11, -1.052619e-11, 
    -1.056695e-11, -1.05553e-11, -1.056722e-11, -1.055964e-11, -1.036891e-11, 
    -1.037838e-11, -1.037326e-11, -1.038288e-11, -1.03761e-11, -1.040622e-11, 
    -1.041525e-11, -1.04575e-11, -1.044017e-11, -1.046775e-11, -1.044297e-11, 
    -1.044736e-11, -1.046865e-11, -1.044431e-11, -1.049754e-11, 
    -1.046145e-11, -1.052849e-11, -1.049245e-11, -1.053075e-11, -1.05238e-11, 
    -1.05353e-11, -1.054561e-11, -1.055858e-11, -1.058249e-11, -1.057696e-11, 
    -1.059696e-11, -1.039249e-11, -1.040476e-11, -1.040368e-11, 
    -1.041652e-11, -1.042602e-11, -1.04466e-11, -1.047961e-11, -1.04672e-11, 
    -1.048998e-11, -1.049455e-11, -1.045994e-11, -1.048119e-11, 
    -1.041297e-11, -1.042399e-11, -1.041743e-11, -1.039345e-11, 
    -1.047005e-11, -1.043075e-11, -1.050332e-11, -1.048204e-11, 
    -1.054414e-11, -1.051326e-11, -1.057391e-11, -1.059982e-11, 
    -1.062421e-11, -1.065269e-11, -1.041146e-11, -1.040312e-11, 
    -1.041805e-11, -1.04387e-11, -1.045787e-11, -1.048333e-11, -1.048594e-11, 
    -1.049071e-11, -1.050307e-11, -1.051345e-11, -1.049221e-11, 
    -1.051606e-11, -1.042654e-11, -1.047346e-11, -1.039997e-11, -1.04221e-11, 
    -1.043749e-11, -1.043074e-11, -1.046578e-11, -1.047404e-11, 
    -1.050758e-11, -1.049024e-11, -1.059342e-11, -1.054778e-11, 
    -1.067438e-11, -1.063902e-11, -1.040021e-11, -1.041143e-11, 
    -1.045048e-11, -1.04319e-11, -1.048503e-11, -1.049811e-11, -1.050874e-11, 
    -1.052231e-11, -1.052378e-11, -1.053183e-11, -1.051864e-11, 
    -1.053131e-11, -1.048339e-11, -1.050481e-11, -1.044602e-11, 
    -1.046033e-11, -1.045375e-11, -1.044653e-11, -1.046882e-11, 
    -1.049255e-11, -1.049306e-11, -1.050067e-11, -1.05221e-11, -1.048525e-11, 
    -1.05993e-11, -1.052887e-11, -1.042367e-11, -1.044528e-11, -1.044837e-11, 
    -1.044e-11, -1.04968e-11, -1.047622e-11, -1.053163e-11, -1.051666e-11, 
    -1.054119e-11, -1.0529e-11, -1.052721e-11, -1.051155e-11, -1.05018e-11, 
    -1.047716e-11, -1.045711e-11, -1.044121e-11, -1.044491e-11, 
    -1.046237e-11, -1.0494e-11, -1.052391e-11, -1.051736e-11, -1.053933e-11, 
    -1.048118e-11, -1.050557e-11, -1.049614e-11, -1.052072e-11, 
    -1.046687e-11, -1.051271e-11, -1.045514e-11, -1.046019e-11, 
    -1.047581e-11, -1.050722e-11, -1.051417e-11, -1.052159e-11, 
    -1.051701e-11, -1.04948e-11, -1.049117e-11, -1.047543e-11, -1.047108e-11, 
    -1.045909e-11, -1.044916e-11, -1.045824e-11, -1.046776e-11, 
    -1.049482e-11, -1.051919e-11, -1.054576e-11, -1.055226e-11, 
    -1.058328e-11, -1.055802e-11, -1.059969e-11, -1.056426e-11, 
    -1.062559e-11, -1.051537e-11, -1.056322e-11, -1.047652e-11, 
    -1.048587e-11, -1.050276e-11, -1.054151e-11, -1.05206e-11, -1.054506e-11, 
    -1.049103e-11, -1.046298e-11, -1.045572e-11, -1.044218e-11, 
    -1.045603e-11, -1.04549e-11, -1.046816e-11, -1.04639e-11, -1.049571e-11, 
    -1.047863e-11, -1.052716e-11, -1.054487e-11, -1.059486e-11, 
    -1.062549e-11, -1.065667e-11, -1.067043e-11, -1.067462e-11, -1.067637e-11 ;

 SMIN_NH4 =
  0.0005315209, 0.0005329163, 0.000532645, 0.0005337701, 0.000533146, 
    0.0005338825, 0.0005318036, 0.0005329712, 0.0005322258, 0.0005316461, 
    0.000535952, 0.0005338199, 0.0005381663, 0.0005368072, 0.0005402206, 
    0.0005379546, 0.0005406773, 0.0005401553, 0.0005417264, 0.0005412763, 
    0.0005432848, 0.000541934, 0.0005443259, 0.0005429623, 0.0005431754, 
    0.0005418892, 0.0005342496, 0.000535687, 0.0005341643, 0.0005343693, 
    0.0005342773, 0.0005331586, 0.0005325946, 0.0005314138, 0.0005316281, 
    0.0005324954, 0.0005344611, 0.0005337939, 0.0005354751, 0.0005354373, 
    0.0005373079, 0.0005364646, 0.0005396078, 0.0005387146, 0.000541295, 
    0.0005406461, 0.0005412644, 0.0005410769, 0.0005412667, 0.0005403151, 
    0.0005407227, 0.0005398854, 0.0005366231, 0.0005375823, 0.0005347204, 
    0.0005329984, 0.0005318546, 0.0005310426, 0.0005311573, 0.0005313761, 
    0.0005325004, 0.0005335573, 0.0005343626, 0.000534901, 0.0005354316, 
    0.0005370368, 0.0005378865, 0.0005397882, 0.0005394452, 0.0005400262, 
    0.0005405815, 0.0005415134, 0.00054136, 0.0005417704, 0.0005400107, 
    0.0005411802, 0.0005392493, 0.0005397775, 0.0005355757, 0.0005339742, 
    0.0005332928, 0.0005326966, 0.0005312455, 0.0005322476, 0.0005318525, 
    0.0005327922, 0.0005333892, 0.0005330939, 0.0005349157, 0.0005342074, 
    0.0005379368, 0.0005363308, 0.0005405168, 0.0005395155, 0.0005407566, 
    0.0005401234, 0.0005412083, 0.0005402318, 0.0005419232, 0.0005422913, 
    0.0005420396, 0.0005430062, 0.0005401773, 0.0005412638, 0.0005330859, 
    0.000533134, 0.0005333584, 0.0005323719, 0.0005323116, 0.0005314076, 
    0.0005322119, 0.0005325543, 0.0005334237, 0.0005339377, 0.0005344262, 
    0.0005355005, 0.0005366997, 0.0005383762, 0.0005395803, 0.0005403872, 
    0.0005398924, 0.0005403291, 0.0005398408, 0.0005396119, 0.0005421532, 
    0.0005407263, 0.0005428671, 0.0005427487, 0.0005417797, 0.0005427618, 
    0.0005331677, 0.0005328906, 0.0005319282, 0.0005326813, 0.000531309, 
    0.0005320771, 0.0005325185, 0.000534222, 0.0005345963, 0.0005349432, 
    0.0005356283, 0.0005365073, 0.0005380489, 0.0005393898, 0.0005406137, 
    0.0005405239, 0.0005405555, 0.0005408286, 0.0005401516, 0.0005409397, 
    0.0005410718, 0.0005407261, 0.0005427326, 0.0005421594, 0.0005427459, 
    0.0005423726, 0.0005329807, 0.0005334468, 0.0005331947, 0.0005336685, 
    0.0005333346, 0.0005348184, 0.000535263, 0.0005373436, 0.0005364899, 
    0.0005378486, 0.0005366279, 0.0005368442, 0.0005378925, 0.0005366938, 
    0.0005393156, 0.000537538, 0.0005408392, 0.0005390645, 0.0005409503, 
    0.0005406079, 0.0005411746, 0.0005416821, 0.0005423204, 0.000543498, 
    0.0005432252, 0.0005442099, 0.0005341417, 0.0005347462, 0.000534693, 
    0.0005353256, 0.0005357932, 0.0005368071, 0.0005384323, 0.0005378211, 
    0.000538943, 0.0005391682, 0.0005374636, 0.0005385101, 0.0005351502, 
    0.000535693, 0.0005353698, 0.0005341885, 0.0005379614, 0.0005360254, 
    0.0005395995, 0.0005385512, 0.0005416095, 0.0005400887, 0.0005430751, 
    0.0005443508, 0.0005455515, 0.0005469536, 0.0005350761, 0.0005346653, 
    0.0005354007, 0.0005364178, 0.0005373615, 0.0005386159, 0.0005387441, 
    0.000538979, 0.0005395874, 0.0005400989, 0.000539053, 0.000540227, 
    0.0005358186, 0.0005381294, 0.0005345092, 0.0005355995, 0.0005363572, 
    0.0005360249, 0.0005377507, 0.0005381572, 0.0005398089, 0.0005389552, 
    0.0005440357, 0.0005417886, 0.0005480213, 0.0005462804, 0.0005345217, 
    0.0005350745, 0.0005369979, 0.0005360829, 0.0005386994, 0.0005393433, 
    0.0005398665, 0.0005405353, 0.0005406074, 0.0005410037, 0.0005403543, 
    0.0005409779, 0.000538618, 0.0005396727, 0.0005367777, 0.0005374823, 
    0.0005371581, 0.0005368023, 0.0005379, 0.0005390688, 0.0005390939, 
    0.0005394685, 0.0005405238, 0.0005387091, 0.000544325, 0.0005408573, 
    0.0005356772, 0.0005367415, 0.0005368936, 0.0005364814, 0.0005392786, 
    0.0005382652, 0.000540994, 0.0005402566, 0.0005414646, 0.0005408644, 
    0.0005407759, 0.0005400049, 0.0005395245, 0.0005383112, 0.0005373236, 
    0.0005365405, 0.0005367225, 0.0005375827, 0.0005391402, 0.0005406133, 
    0.0005402905, 0.0005413721, 0.0005385087, 0.0005397095, 0.0005392453, 
    0.0005404554, 0.0005378047, 0.0005400624, 0.0005372272, 0.0005374759, 
    0.000538245, 0.0005397916, 0.0005401339, 0.0005404991, 0.0005402737, 
    0.0005391802, 0.000539001, 0.0005382259, 0.0005380118, 0.0005374212, 
    0.000536932, 0.0005373788, 0.0005378479, 0.0005391802, 0.0005403804, 
    0.0005416886, 0.0005420087, 0.000543536, 0.0005422924, 0.000544344, 
    0.0005425994, 0.0005456191, 0.0005401933, 0.0005425495, 0.00053828, 
    0.0005387401, 0.0005395722, 0.0005414803, 0.0005404504, 0.0005416548, 
    0.0005389939, 0.0005376124, 0.0005372551, 0.000536588, 0.0005372702, 
    0.0005372147, 0.0005378674, 0.0005376576, 0.0005392243, 0.0005383828, 
    0.0005407729, 0.0005416448, 0.0005441061, 0.000545614, 0.0005471488, 
    0.000547826, 0.0005480321, 0.0005481182 ;

 SMIN_NH4_vr =
  0.002921807, 0.002926611, 0.002925671, 0.002929542, 0.002927392, 
    0.00292992, 0.002922766, 0.002926779, 0.002924214, 0.002922214, 
    0.002937013, 0.00292969, 0.002944614, 0.002939946, 0.002951649, 
    0.002943879, 0.00295321, 0.002951419, 0.002956799, 0.002955253, 
    0.00296212, 0.002957502, 0.002965674, 0.002961013, 0.002961738, 
    0.002957334, 0.002931189, 0.002936124, 0.002930889, 0.002931594, 
    0.002931275, 0.002927423, 0.002925479, 0.002921412, 0.002922146, 
    0.002925131, 0.002931888, 0.002929591, 0.002935367, 0.002935237, 
    0.002941654, 0.00293876, 0.002949539, 0.002946473, 0.002955314, 
    0.002953087, 0.002955203, 0.002954557, 0.002955203, 0.002951944, 
    0.002953334, 0.002950466, 0.002939338, 0.002942626, 0.002932796, 
    0.002926867, 0.002922929, 0.002920134, 0.002920523, 0.002921276, 
    0.002925143, 0.002928776, 0.002931544, 0.00293339, 0.002935209, 
    0.002940719, 0.002943633, 0.00295015, 0.002948974, 0.00295096, 
    0.002952863, 0.002956049, 0.002955523, 0.002956923, 0.002950893, 
    0.002954899, 0.002948278, 0.002950088, 0.002935728, 0.002930224, 
    0.002927877, 0.002925823, 0.002920824, 0.002924274, 0.002922911, 
    0.002926141, 0.002928194, 0.002927174, 0.002933437, 0.002930997, 
    0.002943801, 0.002938289, 0.002952645, 0.002949208, 0.002953458, 
    0.002951289, 0.002954998, 0.002951655, 0.00295744, 0.0029587, 
    0.002957833, 0.002961141, 0.00295145, 0.002955172, 0.002927163, 
    0.002927329, 0.002928097, 0.002924697, 0.002924489, 0.002921373, 
    0.002924138, 0.002925317, 0.002928305, 0.002930068, 0.002931744, 
    0.002935436, 0.00293955, 0.002945299, 0.002949428, 0.002952188, 
    0.002950492, 0.002951984, 0.002950309, 0.00294952, 0.002958219, 
    0.002953334, 0.002960656, 0.002960252, 0.002956932, 0.002960289, 
    0.00292744, 0.002926482, 0.002923168, 0.002925756, 0.002921028, 
    0.002923672, 0.002925187, 0.002931042, 0.002932326, 0.002933519, 
    0.00293587, 0.002938884, 0.002944173, 0.002948767, 0.002952961, 
    0.002952649, 0.002952756, 0.002953687, 0.002951366, 0.002954061, 
    0.002954509, 0.002953326, 0.002960189, 0.002958228, 0.002960231, 
    0.00295895, 0.002926788, 0.002928387, 0.002927516, 0.002929146, 
    0.002927991, 0.002933092, 0.002934616, 0.002941757, 0.002938824, 
    0.002943488, 0.002939292, 0.002940035, 0.002943626, 0.002939511, 
    0.002948503, 0.0029424, 0.00295372, 0.00294763, 0.002954094, 0.002952917, 
    0.002954854, 0.002956592, 0.00295877, 0.002962798, 0.002961859, 
    0.002965227, 0.002930774, 0.002932846, 0.002932663, 0.002934832, 
    0.002936435, 0.002939918, 0.002945491, 0.00294339, 0.002947234, 
    0.002948007, 0.002942154, 0.002945743, 0.002934205, 0.002936064, 
    0.002934954, 0.002930889, 0.002943845, 0.002937194, 0.002949458, 
    0.00294586, 0.002956335, 0.002951126, 0.002961344, 0.002965703, 
    0.002969805, 0.002974583, 0.002933977, 0.002932562, 0.002935085, 
    0.002938577, 0.002941812, 0.002946116, 0.002946553, 0.002947353, 
    0.002949436, 0.002951189, 0.002947599, 0.00295162, 0.002936489, 
    0.002944421, 0.002931985, 0.002935731, 0.002938329, 0.002937189, 
    0.00294311, 0.0029445, 0.002950159, 0.002947234, 0.002964617, 
    0.002956934, 0.00297822, 0.002972281, 0.002932064, 0.00293396, 
    0.002940561, 0.002937421, 0.002946395, 0.002948603, 0.00295039, 
    0.002952681, 0.002952923, 0.00295428, 0.00295205, 0.002954187, 
    0.002946092, 0.002949709, 0.002939774, 0.002942188, 0.002941075, 
    0.002939849, 0.002943612, 0.00294762, 0.002947704, 0.002948982, 
    0.002952592, 0.002946374, 0.002965592, 0.002953724, 0.002936028, 
    0.002939676, 0.002940196, 0.002938782, 0.002948372, 0.002944898, 
    0.002954247, 0.002951717, 0.002955851, 0.002953796, 0.002953486, 
    0.002950846, 0.002949193, 0.002945032, 0.002941637, 0.002938951, 
    0.002939569, 0.002942521, 0.002947856, 0.002952906, 0.002951796, 
    0.002955497, 0.002945681, 0.002949798, 0.002948199, 0.002952348, 
    0.002943321, 0.002951058, 0.002941337, 0.002942186, 0.00294482, 
    0.002950122, 0.002951291, 0.002952542, 0.002951764, 0.002948015, 
    0.002947398, 0.002944736, 0.002943997, 0.002941972, 0.002940286, 
    0.00294182, 0.002943422, 0.002947993, 0.002952102, 0.002956578, 
    0.002957673, 0.002962889, 0.002958635, 0.002965642, 0.002959675, 
    0.002969994, 0.0029515, 0.002959568, 0.002944941, 0.002946515, 
    0.002949364, 0.002955896, 0.002952367, 0.002956491, 0.002947372, 
    0.002942627, 0.002941398, 0.002939109, 0.002941445, 0.002941255, 
    0.002943491, 0.002942767, 0.002948136, 0.002945252, 0.002953436, 
    0.002956422, 0.002964837, 0.002969984, 0.002975223, 0.002977528, 
    0.002978229, 0.00297852,
  0.001884352, 0.00188931, 0.001888347, 0.001892342, 0.001890127, 
    0.001892742, 0.001885358, 0.001889506, 0.001886859, 0.001884799, 
    0.001900082, 0.001892521, 0.001907931, 0.001903118, 0.001915201, 
    0.001907181, 0.001916817, 0.001914972, 0.001920527, 0.001918937, 
    0.001926029, 0.001921261, 0.001929704, 0.001924892, 0.001925644, 
    0.001921103, 0.001894046, 0.001899141, 0.001893743, 0.00189447, 
    0.001894144, 0.001890172, 0.001888168, 0.001883974, 0.001884736, 
    0.001887817, 0.001894797, 0.00189243, 0.001898396, 0.001898262, 
    0.001904893, 0.001901904, 0.001913036, 0.001909876, 0.001919003, 
    0.001916709, 0.001918895, 0.001918233, 0.001918904, 0.001915539, 
    0.001916981, 0.00191402, 0.001902464, 0.001905863, 0.001895717, 
    0.001889602, 0.00188554, 0.001882654, 0.001883062, 0.00188384, 
    0.001887835, 0.00189159, 0.001894449, 0.00189636, 0.001898243, 
    0.00190393, 0.001906942, 0.001913674, 0.001912461, 0.001914516, 
    0.001916481, 0.001919775, 0.001919233, 0.001920684, 0.001914463, 
    0.001918598, 0.00191177, 0.001913639, 0.001898747, 0.001893069, 
    0.001890648, 0.001888532, 0.001883376, 0.001886937, 0.001885533, 
    0.001888873, 0.001890993, 0.001889945, 0.001896412, 0.001893899, 
    0.00190712, 0.00190143, 0.001916252, 0.00191271, 0.001917101, 
    0.001914861, 0.001918697, 0.001915245, 0.001921224, 0.001922524, 
    0.001921635, 0.001925049, 0.001915053, 0.001918894, 0.001889916, 
    0.001890086, 0.001890883, 0.001887379, 0.001887165, 0.001883953, 
    0.001886811, 0.001888028, 0.001891117, 0.001892942, 0.001894676, 
    0.001898487, 0.001902738, 0.001908677, 0.00191294, 0.001915795, 
    0.001914045, 0.00191559, 0.001913862, 0.001913053, 0.001922036, 
    0.001916994, 0.001924558, 0.00192414, 0.001920718, 0.001924188, 
    0.001890207, 0.001889223, 0.001885803, 0.001888479, 0.001883603, 
    0.001886332, 0.001887901, 0.00189395, 0.00189528, 0.00189651, 
    0.001898941, 0.001902057, 0.001907519, 0.001912266, 0.001916596, 
    0.001916279, 0.00191639, 0.001917356, 0.001914962, 0.001917749, 
    0.001918216, 0.001916994, 0.001924084, 0.00192206, 0.001924131, 
    0.001922814, 0.001889543, 0.001891198, 0.001890304, 0.001891985, 
    0.0018908, 0.001896066, 0.001897644, 0.00190502, 0.001901996, 
    0.001906809, 0.001902485, 0.001903252, 0.001906963, 0.00190272, 
    0.001912003, 0.001905709, 0.001917394, 0.001911114, 0.001917787, 
    0.001916577, 0.00191858, 0.001920373, 0.001922629, 0.001926786, 
    0.001925824, 0.001929299, 0.001893666, 0.00189581, 0.001895623, 
    0.001897867, 0.001899525, 0.00190312, 0.001908877, 0.001906713, 
    0.001910686, 0.001911482, 0.001905448, 0.001909153, 0.001897246, 
    0.001899171, 0.001898026, 0.001893834, 0.00190721, 0.00190035, 
    0.00191301, 0.001909301, 0.001920118, 0.00191474, 0.001925294, 
    0.001929794, 0.00193403, 0.001938968, 0.001896982, 0.001895525, 
    0.001898134, 0.001901739, 0.001905085, 0.001909527, 0.001909982, 
    0.001910813, 0.001912966, 0.001914776, 0.001911074, 0.001915229, 
    0.001899614, 0.001907806, 0.001894973, 0.001898839, 0.001901527, 
    0.00190035, 0.001906466, 0.001907906, 0.001913752, 0.001910732, 
    0.001928682, 0.00192075, 0.001942728, 0.001936597, 0.001895015, 
    0.001896977, 0.001903796, 0.001900553, 0.001909824, 0.001912102, 
    0.001913954, 0.001916319, 0.001916575, 0.001917975, 0.00191568, 
    0.001917885, 0.001909536, 0.001913269, 0.001903019, 0.001905515, 
    0.001904367, 0.001903107, 0.001906996, 0.001911132, 0.001911223, 
    0.001912548, 0.001916276, 0.001909861, 0.001929701, 0.001917457, 
    0.001899115, 0.001902887, 0.001903428, 0.001901967, 0.001911874, 
    0.001908287, 0.001917941, 0.001915334, 0.001919605, 0.001917483, 
    0.001917171, 0.001914445, 0.001912746, 0.001908451, 0.001904953, 
    0.001902179, 0.001902824, 0.001905872, 0.001911386, 0.001916597, 
    0.001915456, 0.001919281, 0.001909152, 0.001913401, 0.001911759, 
    0.00191604, 0.001906655, 0.001914642, 0.00190461, 0.001905492, 
    0.001908215, 0.001913688, 0.001914901, 0.001916192, 0.001915396, 
    0.001911526, 0.001910893, 0.00190815, 0.001907391, 0.0019053, 
    0.001903567, 0.00190515, 0.001906811, 0.001911529, 0.001915774, 
    0.001920398, 0.00192153, 0.00192692, 0.00192253, 0.001929769, 
    0.001923611, 0.001934267, 0.001915108, 0.001923434, 0.00190834, 
    0.001909969, 0.001912912, 0.001919659, 0.00191602, 0.001920277, 
    0.001910868, 0.001905976, 0.001904711, 0.001902347, 0.001904765, 
    0.001904569, 0.001906881, 0.001906138, 0.001911685, 0.001908707, 
    0.001917163, 0.001920243, 0.001928934, 0.001934251, 0.001939659, 
    0.001942043, 0.001942768, 0.001943072,
  0.001890095, 0.001895119, 0.001894143, 0.001898192, 0.001895947, 
    0.001898597, 0.001891115, 0.001895318, 0.001892635, 0.001890548, 
    0.001906039, 0.001898373, 0.001913996, 0.001909114, 0.00192137, 
    0.001913236, 0.001923009, 0.001921137, 0.001926772, 0.001925158, 
    0.001932357, 0.001927517, 0.001936086, 0.001931202, 0.001931966, 
    0.001927357, 0.001899918, 0.001905084, 0.001899611, 0.001900348, 
    0.001900018, 0.001895993, 0.001893962, 0.001889712, 0.001890484, 
    0.001893606, 0.00190068, 0.00189828, 0.001904328, 0.001904191, 
    0.001910914, 0.001907884, 0.001919173, 0.001915967, 0.001925226, 
    0.001922899, 0.001925116, 0.001924444, 0.001925125, 0.001921712, 
    0.001923174, 0.00192017, 0.001908451, 0.001911898, 0.001901612, 
    0.001895415, 0.001891299, 0.001888375, 0.001888788, 0.001889576, 
    0.001893625, 0.001897429, 0.001900326, 0.001902263, 0.001904172, 
    0.001909939, 0.001912992, 0.00191982, 0.00191859, 0.001920674, 
    0.001922667, 0.001926009, 0.00192546, 0.001926931, 0.00192062, 
    0.001924815, 0.001917888, 0.001919784, 0.001904686, 0.001898928, 
    0.001896475, 0.001894331, 0.001889106, 0.001892714, 0.001891292, 
    0.001894676, 0.001896824, 0.001895762, 0.001902316, 0.001899769, 
    0.001913173, 0.001907404, 0.001922435, 0.001918842, 0.001923296, 
    0.001921024, 0.001924915, 0.001921413, 0.001927479, 0.001928799, 
    0.001927897, 0.001931361, 0.001921219, 0.001925116, 0.001895732, 
    0.001895905, 0.001896713, 0.001893162, 0.001892945, 0.00188969, 
    0.001892587, 0.00189382, 0.001896949, 0.001898799, 0.001900556, 
    0.001904419, 0.00190873, 0.001914752, 0.001919075, 0.001921971, 
    0.001920196, 0.001921763, 0.001920011, 0.001919189, 0.001928304, 
    0.001923188, 0.001930863, 0.001930439, 0.001926966, 0.001930487, 
    0.001896027, 0.00189503, 0.001891565, 0.001894277, 0.001889336, 
    0.001892102, 0.001893691, 0.001899821, 0.001901168, 0.001902416, 
    0.001904879, 0.001908039, 0.001913577, 0.001918392, 0.001922783, 
    0.001922462, 0.001922575, 0.001923555, 0.001921126, 0.001923954, 
    0.001924428, 0.001923188, 0.001930382, 0.001928328, 0.00193043, 
    0.001929093, 0.001895354, 0.001897032, 0.001896125, 0.00189783, 
    0.001896629, 0.001901966, 0.001903565, 0.001911043, 0.001907977, 
    0.001912858, 0.001908473, 0.00190925, 0.001913015, 0.00190871, 
    0.001918125, 0.001911743, 0.001923593, 0.001917224, 0.001923992, 
    0.001922764, 0.001924797, 0.001926616, 0.001928905, 0.001933124, 
    0.001932148, 0.001935675, 0.001899533, 0.001901707, 0.001901516, 
    0.001903791, 0.001905472, 0.001909116, 0.001914954, 0.00191276, 
    0.001916788, 0.001917596, 0.001911476, 0.001915234, 0.001903162, 
    0.001905113, 0.001903952, 0.001899704, 0.001913264, 0.001906309, 
    0.001919146, 0.001915384, 0.001926357, 0.001920902, 0.00193161, 
    0.001936178, 0.001940478, 0.001945493, 0.001902894, 0.001901417, 
    0.001904062, 0.001907717, 0.001911109, 0.001915613, 0.001916074, 
    0.001916918, 0.001919102, 0.001920937, 0.001917183, 0.001921397, 
    0.001905564, 0.001913868, 0.001900858, 0.001904777, 0.001907502, 
    0.001906308, 0.001912509, 0.00191397, 0.001919899, 0.001916835, 
    0.00193505, 0.001926999, 0.001949312, 0.001943086, 0.001900901, 
    0.001902889, 0.001909802, 0.001906514, 0.001915914, 0.001918225, 
    0.001920104, 0.001922503, 0.001922762, 0.001924183, 0.001921854, 
    0.001924091, 0.001915623, 0.001919409, 0.001909013, 0.001911545, 
    0.001910381, 0.001909103, 0.001913046, 0.001917242, 0.001917333, 
    0.001918678, 0.001922462, 0.001915952, 0.001936086, 0.001923659, 
    0.001905056, 0.001908881, 0.001909428, 0.001907947, 0.001917993, 
    0.001914355, 0.001924149, 0.001921504, 0.001925837, 0.001923684, 
    0.001923367, 0.001920601, 0.001918878, 0.001914522, 0.001910975, 
    0.001908162, 0.001908817, 0.001911907, 0.001917499, 0.001922785, 
    0.001921627, 0.001925508, 0.001915233, 0.001919543, 0.001917877, 
    0.00192222, 0.001912701, 0.001920804, 0.001910627, 0.001911521, 
    0.001914283, 0.001919835, 0.001921064, 0.001922374, 0.001921566, 
    0.001917641, 0.001916999, 0.001914216, 0.001913447, 0.001911327, 
    0.001909569, 0.001911175, 0.001912859, 0.001917643, 0.00192195, 
    0.001926642, 0.00192779, 0.001933262, 0.001928806, 0.001936155, 
    0.001929905, 0.00194072, 0.001921275, 0.001929724, 0.001914409, 
    0.001916062, 0.001919048, 0.001925892, 0.0019222, 0.001926519, 
    0.001916974, 0.001912012, 0.00191073, 0.001908333, 0.001910784, 
    0.001910585, 0.00191293, 0.001912177, 0.001917802, 0.001914781, 
    0.001923359, 0.001926485, 0.001935305, 0.001940703, 0.001946194, 
    0.001948616, 0.001949352, 0.00194966,
  0.001831809, 0.001836763, 0.0018358, 0.001839794, 0.001837579, 0.001840193, 
    0.001832814, 0.001836959, 0.001834313, 0.001832255, 0.001847539, 
    0.001839972, 0.001855395, 0.001850573, 0.001862682, 0.001854645, 
    0.001864302, 0.001862451, 0.001868022, 0.001866426, 0.001873548, 
    0.001868759, 0.001877238, 0.001872405, 0.001873161, 0.0018686, 
    0.001841496, 0.001846597, 0.001841193, 0.001841921, 0.001841595, 
    0.001837624, 0.001835622, 0.001831431, 0.001832192, 0.001835271, 
    0.001842248, 0.001839881, 0.001845847, 0.001845713, 0.001852351, 
    0.001849358, 0.001860509, 0.001857341, 0.001866493, 0.001864192, 
    0.001866385, 0.00186572, 0.001866394, 0.001863019, 0.001864465, 
    0.001861495, 0.001849919, 0.001853322, 0.001843168, 0.001837056, 
    0.001832995, 0.001830113, 0.00183052, 0.001831297, 0.001835289, 
    0.001839041, 0.001841899, 0.00184381, 0.001845693, 0.001851389, 
    0.001854404, 0.001861149, 0.001859933, 0.001861994, 0.001863963, 
    0.001867268, 0.001866724, 0.00186818, 0.00186194, 0.001866087, 
    0.00185924, 0.001861113, 0.001846203, 0.001840519, 0.001838101, 
    0.001835985, 0.001830834, 0.001834391, 0.001832989, 0.001836325, 
    0.001838444, 0.001837396, 0.001843863, 0.001841349, 0.001854582, 
    0.001848885, 0.001863734, 0.001860183, 0.001864585, 0.001862339, 
    0.001866187, 0.001862724, 0.001868722, 0.001870027, 0.001869135, 
    0.001872562, 0.001862532, 0.001866385, 0.001837367, 0.001837538, 
    0.001838334, 0.001834833, 0.001834619, 0.00183141, 0.001834265, 
    0.001835481, 0.001838567, 0.001840392, 0.001842126, 0.001845938, 
    0.001850194, 0.001856142, 0.001860413, 0.001863275, 0.00186152, 
    0.001863069, 0.001861337, 0.001860526, 0.001869538, 0.001864478, 
    0.001872069, 0.001871649, 0.001868215, 0.001871697, 0.001837658, 
    0.001836674, 0.001833258, 0.001835932, 0.00183106, 0.001833787, 
    0.001835354, 0.001841401, 0.00184273, 0.001843961, 0.001846392, 
    0.001849512, 0.001854981, 0.001859738, 0.001864078, 0.00186376, 
    0.001863872, 0.001864841, 0.00186244, 0.001865235, 0.001865704, 
    0.001864478, 0.001871593, 0.001869561, 0.00187164, 0.001870317, 
    0.001836994, 0.001838649, 0.001837755, 0.001839436, 0.001838251, 
    0.001843518, 0.001845096, 0.001852479, 0.00184945, 0.00185427, 
    0.00184994, 0.001850707, 0.001854427, 0.001850174, 0.001859475, 
    0.00185317, 0.001864879, 0.001858585, 0.001865273, 0.001864059, 
    0.001866069, 0.001867868, 0.001870132, 0.001874307, 0.00187334, 
    0.001876831, 0.001841116, 0.001843261, 0.001843073, 0.001845318, 
    0.001846978, 0.001850575, 0.001856341, 0.001854173, 0.001858153, 
    0.001858952, 0.001852905, 0.001856618, 0.001844697, 0.001846624, 
    0.001845477, 0.001841285, 0.001854672, 0.001847804, 0.001860483, 
    0.001856766, 0.001867612, 0.001862219, 0.001872808, 0.00187733, 
    0.001881586, 0.001886555, 0.001844432, 0.001842975, 0.001845585, 
    0.001849194, 0.001852543, 0.001856992, 0.001857448, 0.001858281, 
    0.001860439, 0.001862253, 0.001858544, 0.001862708, 0.00184707, 
    0.001855268, 0.001842423, 0.001846293, 0.001848981, 0.001847802, 
    0.001853926, 0.001855368, 0.001861227, 0.001858199, 0.001876214, 
    0.001868248, 0.001890338, 0.00188417, 0.001842465, 0.001844428, 
    0.001851253, 0.001848006, 0.001857289, 0.001859573, 0.001861429, 
    0.001863801, 0.001864057, 0.001865462, 0.00186316, 0.001865371, 
    0.001857002, 0.001860743, 0.001850473, 0.001852974, 0.001851824, 
    0.001850562, 0.001854456, 0.001858602, 0.001858691, 0.00186002, 
    0.001863763, 0.001857327, 0.001877241, 0.001864947, 0.001846567, 
    0.001850343, 0.001850883, 0.00184942, 0.001859344, 0.00185575, 
    0.001865428, 0.001862813, 0.001867097, 0.001864969, 0.001864655, 
    0.001861921, 0.001860218, 0.001855914, 0.001852411, 0.001849633, 
    0.001850279, 0.001853331, 0.001858856, 0.00186408, 0.001862936, 
    0.001866772, 0.001856617, 0.001860876, 0.00185923, 0.001863522, 
    0.001854116, 0.001862124, 0.001852067, 0.001852949, 0.001855678, 
    0.001861164, 0.001862379, 0.001863674, 0.001862875, 0.001858996, 
    0.001858361, 0.001855612, 0.001854853, 0.001852758, 0.001851022, 
    0.001852607, 0.001854272, 0.001858998, 0.001863255, 0.001867894, 
    0.001869029, 0.001874444, 0.001870036, 0.001877309, 0.001871125, 
    0.001881828, 0.001862589, 0.001870944, 0.001855802, 0.001857435, 
    0.001860386, 0.001867153, 0.001863501, 0.001867773, 0.001858336, 
    0.001853436, 0.001852168, 0.001849802, 0.001852222, 0.001852025, 
    0.001854341, 0.001853597, 0.001859155, 0.00185617, 0.001864647, 
    0.001867739, 0.001876465, 0.00188181, 0.001887248, 0.001889648, 
    0.001890378, 0.001890683,
  0.001659499, 0.001664149, 0.001663245, 0.001666996, 0.001664915, 
    0.001667371, 0.001660441, 0.001664333, 0.001661849, 0.001659917, 
    0.001674279, 0.001667163, 0.001681673, 0.001677133, 0.001688542, 
    0.001680967, 0.00169007, 0.001688323, 0.001693581, 0.001692075, 
    0.001698802, 0.001694276, 0.00170229, 0.001697721, 0.001698436, 
    0.001694127, 0.001668595, 0.001673393, 0.001668311, 0.001668995, 
    0.001668688, 0.001664958, 0.001663079, 0.001659143, 0.001659858, 
    0.001662748, 0.001669302, 0.001667077, 0.001672686, 0.001672559, 
    0.001678806, 0.001675989, 0.001686493, 0.001683507, 0.001692137, 
    0.001689966, 0.001692035, 0.001691408, 0.001692044, 0.00168886, 
    0.001690224, 0.001687422, 0.001676516, 0.001679721, 0.001670166, 
    0.001664425, 0.001660612, 0.001657907, 0.001658289, 0.001659018, 
    0.001662765, 0.001666288, 0.001668974, 0.00167077, 0.001672541, 
    0.001677902, 0.00168074, 0.001687097, 0.001685949, 0.001687893, 
    0.00168975, 0.001692869, 0.001692356, 0.00169373, 0.001687842, 
    0.001691755, 0.001685295, 0.001687062, 0.001673023, 0.001667677, 
    0.001665406, 0.001663418, 0.001658584, 0.001661922, 0.001660606, 
    0.001663737, 0.001665728, 0.001664743, 0.001670819, 0.001668457, 
    0.001680908, 0.001675543, 0.001689534, 0.001686185, 0.001690337, 
    0.001688218, 0.001691848, 0.001688581, 0.001694242, 0.001695475, 
    0.001694632, 0.001697869, 0.0016884, 0.001692035, 0.001664716, 
    0.001664876, 0.001665624, 0.001662337, 0.001662136, 0.001659124, 
    0.001661804, 0.001662945, 0.001665843, 0.001667557, 0.001669187, 
    0.001672771, 0.001676776, 0.001682376, 0.001686402, 0.001689101, 
    0.001687446, 0.001688907, 0.001687273, 0.001686508, 0.001695013, 
    0.001690237, 0.001697403, 0.001697007, 0.001693763, 0.001697051, 
    0.001664989, 0.001664065, 0.001660858, 0.001663368, 0.001658796, 
    0.001661355, 0.001662827, 0.001668506, 0.001669755, 0.001670912, 
    0.001673198, 0.001676133, 0.001681283, 0.001685765, 0.001689858, 
    0.001689558, 0.001689664, 0.001690579, 0.001688313, 0.00169095, 
    0.001691393, 0.001690236, 0.001696954, 0.001695034, 0.001696998, 
    0.001695748, 0.001664365, 0.00166592, 0.00166508, 0.00166666, 
    0.001665547, 0.001670496, 0.00167198, 0.001678927, 0.001676075, 
    0.001680614, 0.001676536, 0.001677259, 0.001680762, 0.001676757, 
    0.001685518, 0.001679578, 0.001690614, 0.00168468, 0.001690986, 
    0.001689841, 0.001691737, 0.001693436, 0.001695573, 0.001699518, 
    0.001698605, 0.001701905, 0.001668238, 0.001670255, 0.001670077, 
    0.001672188, 0.001673749, 0.001677134, 0.001682564, 0.001680522, 
    0.001684271, 0.001685024, 0.001679328, 0.001682825, 0.001671604, 
    0.001673417, 0.001672338, 0.001668397, 0.001680992, 0.001674527, 
    0.001686468, 0.001682964, 0.001693194, 0.001688105, 0.001698102, 
    0.001702378, 0.001706403, 0.00171111, 0.001671355, 0.001669985, 
    0.001672439, 0.001675835, 0.001678986, 0.001683178, 0.001683606, 
    0.001684392, 0.001686426, 0.001688137, 0.00168464, 0.001688566, 
    0.001673837, 0.001681554, 0.001669467, 0.001673105, 0.001675635, 
    0.001674525, 0.001680288, 0.001681647, 0.00168717, 0.001684315, 
    0.001701323, 0.001693795, 0.001714694, 0.00170885, 0.001669506, 
    0.001671351, 0.001677772, 0.001674716, 0.001683457, 0.00168561, 
    0.00168736, 0.001689597, 0.001689839, 0.001691165, 0.001688992, 
    0.001691079, 0.001683187, 0.001686713, 0.001677038, 0.001679392, 
    0.001678309, 0.001677121, 0.001680788, 0.001684695, 0.001684779, 
    0.001686032, 0.001689564, 0.001683493, 0.001702294, 0.00169068, 
    0.001673362, 0.001676916, 0.001677424, 0.001676047, 0.001685394, 
    0.001682007, 0.001691132, 0.001688665, 0.001692708, 0.001690699, 
    0.001690403, 0.001687824, 0.001686218, 0.001682162, 0.001678863, 
    0.001676247, 0.001676855, 0.001679729, 0.001684934, 0.001689861, 
    0.001688781, 0.0016924, 0.001682824, 0.001686838, 0.001685287, 
    0.001689333, 0.001680468, 0.001688017, 0.001678538, 0.001679369, 
    0.001681939, 0.001687111, 0.001688255, 0.001689477, 0.001688723, 
    0.001685066, 0.001684467, 0.001681877, 0.001681162, 0.001679188, 
    0.001677555, 0.001679047, 0.001680615, 0.001685068, 0.001689082, 
    0.00169346, 0.001694532, 0.00169965, 0.001695483, 0.001702359, 
    0.001696514, 0.001706635, 0.001688455, 0.001696341, 0.001682056, 
    0.001683595, 0.001686377, 0.001692762, 0.001689314, 0.001693346, 
    0.001684444, 0.001679828, 0.001678634, 0.001676406, 0.001678684, 
    0.001678499, 0.00168068, 0.001679979, 0.001685216, 0.001682403, 
    0.001690396, 0.001693314, 0.001701559, 0.001706616, 0.001711765, 
    0.00171404, 0.001714732, 0.001715021,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.822918e-06, 1.832765e-06, 1.830849e-06, 1.838805e-06, 1.83439e-06, 
    1.839602e-06, 1.824912e-06, 1.833155e-06, 1.827891e-06, 1.823803e-06, 
    1.854285e-06, 1.839159e-06, 1.870063e-06, 1.860371e-06, 1.884762e-06, 
    1.868552e-06, 1.888038e-06, 1.884294e-06, 1.895575e-06, 1.89234e-06, 
    1.906798e-06, 1.897068e-06, 1.914314e-06, 1.904473e-06, 1.90601e-06, 
    1.896746e-06, 1.842201e-06, 1.8524e-06, 1.841597e-06, 1.84305e-06, 
    1.842398e-06, 1.83448e-06, 1.830495e-06, 1.822166e-06, 1.823677e-06, 
    1.829795e-06, 1.843702e-06, 1.838976e-06, 1.850898e-06, 1.850629e-06, 
    1.86394e-06, 1.857933e-06, 1.880372e-06, 1.873982e-06, 1.892474e-06, 
    1.887816e-06, 1.892255e-06, 1.890908e-06, 1.892272e-06, 1.885442e-06, 
    1.888367e-06, 1.882362e-06, 1.859059e-06, 1.865894e-06, 1.84554e-06, 
    1.833347e-06, 1.825273e-06, 1.819552e-06, 1.82036e-06, 1.821901e-06, 
    1.829831e-06, 1.837302e-06, 1.843004e-06, 1.846823e-06, 1.850589e-06, 
    1.862008e-06, 1.868067e-06, 1.881664e-06, 1.879208e-06, 1.88337e-06, 
    1.887352e-06, 1.894045e-06, 1.892942e-06, 1.895893e-06, 1.883261e-06, 
    1.891651e-06, 1.877808e-06, 1.88159e-06, 1.851611e-06, 1.840252e-06, 
    1.835429e-06, 1.831216e-06, 1.820981e-06, 1.828046e-06, 1.825259e-06, 
    1.831892e-06, 1.836113e-06, 1.834025e-06, 1.846927e-06, 1.841906e-06, 
    1.868426e-06, 1.856982e-06, 1.886888e-06, 1.879712e-06, 1.888609e-06, 
    1.884067e-06, 1.891853e-06, 1.884845e-06, 1.896992e-06, 1.899641e-06, 
    1.89783e-06, 1.904791e-06, 1.884456e-06, 1.892253e-06, 1.833967e-06, 
    1.834307e-06, 1.835894e-06, 1.828924e-06, 1.828498e-06, 1.822123e-06, 
    1.827795e-06, 1.830212e-06, 1.836357e-06, 1.839995e-06, 1.843457e-06, 
    1.851079e-06, 1.859608e-06, 1.871564e-06, 1.880177e-06, 1.885959e-06, 
    1.882412e-06, 1.885543e-06, 1.882043e-06, 1.880404e-06, 1.898647e-06, 
    1.888393e-06, 1.903789e-06, 1.902936e-06, 1.895962e-06, 1.903031e-06, 
    1.834546e-06, 1.832587e-06, 1.825793e-06, 1.831109e-06, 1.821429e-06, 
    1.826844e-06, 1.82996e-06, 1.84201e-06, 1.844663e-06, 1.847123e-06, 
    1.851988e-06, 1.858239e-06, 1.869228e-06, 1.878813e-06, 1.887584e-06, 
    1.88694e-06, 1.887167e-06, 1.889128e-06, 1.884271e-06, 1.889925e-06, 
    1.890874e-06, 1.888392e-06, 1.902821e-06, 1.898694e-06, 1.902917e-06, 
    1.900229e-06, 1.833224e-06, 1.83652e-06, 1.834738e-06, 1.838089e-06, 
    1.835728e-06, 1.846237e-06, 1.849394e-06, 1.864196e-06, 1.858115e-06, 
    1.867798e-06, 1.859098e-06, 1.860638e-06, 1.868112e-06, 1.859568e-06, 
    1.878283e-06, 1.865583e-06, 1.889204e-06, 1.876487e-06, 1.890001e-06, 
    1.887545e-06, 1.891613e-06, 1.89526e-06, 1.899853e-06, 1.90834e-06, 
    1.906373e-06, 1.913481e-06, 1.84144e-06, 1.845725e-06, 1.845348e-06, 
    1.849837e-06, 1.85316e-06, 1.860372e-06, 1.871966e-06, 1.867603e-06, 
    1.875617e-06, 1.877227e-06, 1.865053e-06, 1.872523e-06, 1.848594e-06, 
    1.85245e-06, 1.850154e-06, 1.841776e-06, 1.868605e-06, 1.854813e-06, 
    1.880317e-06, 1.872819e-06, 1.894739e-06, 1.883823e-06, 1.90529e-06, 
    1.914499e-06, 1.923188e-06, 1.93336e-06, 1.848066e-06, 1.845152e-06, 
    1.850371e-06, 1.857602e-06, 1.864324e-06, 1.873277e-06, 1.874195e-06, 
    1.875874e-06, 1.880229e-06, 1.883893e-06, 1.876404e-06, 1.884812e-06, 
    1.853343e-06, 1.869805e-06, 1.844048e-06, 1.851786e-06, 1.857174e-06, 
    1.85481e-06, 1.867102e-06, 1.870004e-06, 1.881818e-06, 1.875707e-06, 
    1.912223e-06, 1.896028e-06, 1.941124e-06, 1.928473e-06, 1.844134e-06, 
    1.848056e-06, 1.861733e-06, 1.85522e-06, 1.873876e-06, 1.878481e-06, 
    1.882228e-06, 1.887022e-06, 1.887541e-06, 1.890385e-06, 1.885725e-06, 
    1.8902e-06, 1.873295e-06, 1.880841e-06, 1.860167e-06, 1.865189e-06, 
    1.862878e-06, 1.860344e-06, 1.868169e-06, 1.87652e-06, 1.8767e-06, 
    1.879381e-06, 1.886944e-06, 1.873949e-06, 1.914315e-06, 1.889338e-06, 
    1.852336e-06, 1.859907e-06, 1.860991e-06, 1.858055e-06, 1.878018e-06, 
    1.870774e-06, 1.890315e-06, 1.885025e-06, 1.893696e-06, 1.889385e-06, 
    1.888751e-06, 1.883221e-06, 1.879781e-06, 1.871104e-06, 1.864057e-06, 
    1.858479e-06, 1.859776e-06, 1.865906e-06, 1.877031e-06, 1.887585e-06, 
    1.885271e-06, 1.893035e-06, 1.872517e-06, 1.881108e-06, 1.877785e-06, 
    1.886454e-06, 1.867486e-06, 1.883632e-06, 1.863368e-06, 1.865141e-06, 
    1.87063e-06, 1.881692e-06, 1.884145e-06, 1.886764e-06, 1.885148e-06, 
    1.877316e-06, 1.876034e-06, 1.870495e-06, 1.868967e-06, 1.864754e-06, 
    1.861267e-06, 1.864452e-06, 1.867798e-06, 1.877318e-06, 1.885916e-06, 
    1.89531e-06, 1.897612e-06, 1.908618e-06, 1.899655e-06, 1.914453e-06, 
    1.901866e-06, 1.923681e-06, 1.884571e-06, 1.901501e-06, 1.87088e-06, 
    1.874168e-06, 1.880121e-06, 1.89381e-06, 1.886415e-06, 1.895065e-06, 
    1.875984e-06, 1.866117e-06, 1.863569e-06, 1.858818e-06, 1.863678e-06, 
    1.863282e-06, 1.867937e-06, 1.866441e-06, 1.877634e-06, 1.871618e-06, 
    1.888732e-06, 1.894995e-06, 1.912734e-06, 1.923643e-06, 1.93478e-06, 
    1.939705e-06, 1.941205e-06, 1.941833e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.069113e-06, 8.103319e-06, 8.096653e-06, 8.124252e-06, 8.108936e-06, 
    8.126992e-06, 8.076011e-06, 8.104614e-06, 8.086345e-06, 8.07213e-06, 
    8.177773e-06, 8.125418e-06, 8.232298e-06, 8.198826e-06, 8.282937e-06, 
    8.227056e-06, 8.294209e-06, 8.281319e-06, 8.320124e-06, 8.308991e-06, 
    8.358618e-06, 8.325235e-06, 8.384383e-06, 8.350637e-06, 8.355897e-06, 
    8.32409e-06, 8.136024e-06, 8.171308e-06, 8.133915e-06, 8.138946e-06, 
    8.136682e-06, 8.10921e-06, 8.095366e-06, 8.066435e-06, 8.071675e-06, 
    8.092924e-06, 8.141147e-06, 8.124765e-06, 8.166056e-06, 8.165125e-06, 
    8.211126e-06, 8.190372e-06, 8.267803e-06, 8.245768e-06, 8.309446e-06, 
    8.293406e-06, 8.308672e-06, 8.30403e-06, 8.308708e-06, 8.285208e-06, 
    8.295257e-06, 8.27459e-06, 8.194354e-06, 8.217955e-06, 8.147559e-06, 
    8.105258e-06, 8.077227e-06, 8.057345e-06, 8.060138e-06, 8.065494e-06, 
    8.093031e-06, 8.118953e-06, 8.138721e-06, 8.151936e-06, 8.164966e-06, 
    8.204423e-06, 8.225351e-06, 8.272229e-06, 8.263773e-06, 8.278091e-06, 
    8.291802e-06, 8.314806e-06, 8.311015e-06, 8.321143e-06, 8.277679e-06, 
    8.306549e-06, 8.258882e-06, 8.271909e-06, 8.168538e-06, 8.129222e-06, 
    8.112474e-06, 8.097856e-06, 8.062291e-06, 8.086839e-06, 8.077149e-06, 
    8.10018e-06, 8.114818e-06, 8.107565e-06, 8.152289e-06, 8.134878e-06, 
    8.226579e-06, 8.187051e-06, 8.290213e-06, 8.265491e-06, 8.296116e-06, 
    8.280485e-06, 8.307251e-06, 8.283147e-06, 8.324904e-06, 8.334002e-06, 
    8.327766e-06, 8.351675e-06, 8.281756e-06, 8.308582e-06, 8.107409e-06, 
    8.108591e-06, 8.114086e-06, 8.089874e-06, 8.088394e-06, 8.066238e-06, 
    8.085934e-06, 8.094327e-06, 8.115649e-06, 8.128249e-06, 8.140236e-06, 
    8.166632e-06, 8.19611e-06, 8.237387e-06, 8.267081e-06, 8.286985e-06, 
    8.274772e-06, 8.285538e-06, 8.273482e-06, 8.267824e-06, 8.330565e-06, 
    8.295315e-06, 8.348211e-06, 8.345285e-06, 8.321315e-06, 8.345591e-06, 
    8.109404e-06, 8.102597e-06, 8.078997e-06, 8.09745e-06, 8.06381e-06, 
    8.082625e-06, 8.093431e-06, 8.135217e-06, 8.14441e-06, 8.152931e-06, 
    8.169763e-06, 8.191369e-06, 8.229316e-06, 8.262362e-06, 8.292568e-06, 
    8.290343e-06, 8.291117e-06, 8.297849e-06, 8.281131e-06, 8.300578e-06, 
    8.303828e-06, 8.295295e-06, 8.344868e-06, 8.330697e-06, 8.345189e-06, 
    8.335948e-06, 8.104797e-06, 8.11622e-06, 8.110028e-06, 8.12165e-06, 
    8.11344e-06, 8.149864e-06, 8.160779e-06, 8.21195e-06, 8.190939e-06, 
    8.224385e-06, 8.194323e-06, 8.199643e-06, 8.225424e-06, 8.195927e-06, 
    8.260501e-06, 8.216674e-06, 8.298101e-06, 8.254272e-06, 8.300831e-06, 
    8.292368e-06, 8.306353e-06, 8.318889e-06, 8.334653e-06, 8.363776e-06, 
    8.357015e-06, 8.38139e-06, 8.133271e-06, 8.148097e-06, 8.146797e-06, 
    8.162327e-06, 8.173812e-06, 8.198757e-06, 8.238772e-06, 8.223707e-06, 
    8.251346e-06, 8.256898e-06, 8.21488e-06, 8.240652e-06, 8.157953e-06, 
    8.171276e-06, 8.16334e-06, 8.134305e-06, 8.22709e-06, 8.179422e-06, 
    8.267469e-06, 8.24161e-06, 8.317075e-06, 8.279513e-06, 8.353295e-06, 
    8.384854e-06, 8.414617e-06, 8.44936e-06, 8.1562e-06, 8.1461e-06, 
    8.164162e-06, 8.189162e-06, 8.212384e-06, 8.243286e-06, 8.246444e-06, 
    8.252219e-06, 8.26722e-06, 8.279841e-06, 8.254019e-06, 8.282983e-06, 
    8.174337e-06, 8.231231e-06, 8.142167e-06, 8.168948e-06, 8.187574e-06, 
    8.179407e-06, 8.22188e-06, 8.231882e-06, 8.272591e-06, 8.251544e-06, 
    8.377029e-06, 8.321458e-06, 8.475862e-06, 8.43265e-06, 8.142564e-06, 
    8.156135e-06, 8.203421e-06, 8.180914e-06, 8.245331e-06, 8.261204e-06, 
    8.274102e-06, 8.290603e-06, 8.292373e-06, 8.302156e-06, 8.286111e-06, 
    8.30151e-06, 8.243261e-06, 8.269276e-06, 8.197932e-06, 8.215264e-06, 
    8.207284e-06, 8.198515e-06, 8.225531e-06, 8.254327e-06, 8.254949e-06, 
    8.26417e-06, 8.290166e-06, 8.245436e-06, 8.384141e-06, 8.298381e-06, 
    8.170942e-06, 8.197093e-06, 8.200842e-06, 8.190702e-06, 8.259588e-06, 
    8.234608e-06, 8.301919e-06, 8.283704e-06, 8.313526e-06, 8.298699e-06, 
    8.296498e-06, 8.277468e-06, 8.2656e-06, 8.235682e-06, 8.21134e-06, 
    8.192074e-06, 8.196536e-06, 8.217708e-06, 8.256068e-06, 8.292423e-06, 
    8.284444e-06, 8.311151e-06, 8.240481e-06, 8.270088e-06, 8.258618e-06, 
    8.288487e-06, 8.223268e-06, 8.278898e-06, 8.209045e-06, 8.215156e-06, 
    8.234088e-06, 8.272214e-06, 8.28066e-06, 8.289671e-06, 8.284097e-06, 
    8.25711e-06, 8.252686e-06, 8.233575e-06, 8.228284e-06, 8.213748e-06, 
    8.201687e-06, 8.212687e-06, 8.224216e-06, 8.257061e-06, 8.28666e-06, 
    8.31896e-06, 8.326874e-06, 8.364607e-06, 8.333849e-06, 8.384573e-06, 
    8.341392e-06, 8.416167e-06, 8.282125e-06, 8.340334e-06, 8.234957e-06, 
    8.246287e-06, 8.266788e-06, 8.313881e-06, 8.288451e-06, 8.31819e-06, 
    8.252508e-06, 8.218443e-06, 8.209648e-06, 8.19323e-06, 8.210006e-06, 
    8.208643e-06, 8.224709e-06, 8.21953e-06, 8.258127e-06, 8.237386e-06, 
    8.296326e-06, 8.317858e-06, 8.378731e-06, 8.41607e-06, 8.45415e-06, 
    8.470949e-06, 8.476066e-06, 8.478196e-06,
  5.553977e-06, 5.583309e-06, 5.577607e-06, 5.601284e-06, 5.588151e-06, 
    5.603656e-06, 5.559926e-06, 5.58447e-06, 5.568801e-06, 5.556623e-06, 
    5.647299e-06, 5.602342e-06, 5.694154e-06, 5.665396e-06, 5.737729e-06, 
    5.68967e-06, 5.747435e-06, 5.736354e-06, 5.769754e-06, 5.760181e-06, 
    5.802933e-06, 5.774174e-06, 5.825147e-06, 5.796068e-06, 5.80061e-06, 
    5.773224e-06, 5.611393e-06, 5.641692e-06, 5.609596e-06, 5.613914e-06, 
    5.611979e-06, 5.588417e-06, 5.576547e-06, 5.551745e-06, 5.556248e-06, 
    5.574469e-06, 5.615857e-06, 5.601806e-06, 5.63726e-06, 5.636459e-06, 
    5.675994e-06, 5.658159e-06, 5.724733e-06, 5.705793e-06, 5.760581e-06, 
    5.746787e-06, 5.75993e-06, 5.755945e-06, 5.759982e-06, 5.739756e-06, 
    5.748419e-06, 5.730634e-06, 5.661496e-06, 5.681788e-06, 5.621322e-06, 
    5.585035e-06, 5.560999e-06, 5.543953e-06, 5.546362e-06, 5.550952e-06, 
    5.574576e-06, 5.596823e-06, 5.61379e-06, 5.625146e-06, 5.636344e-06, 
    5.670244e-06, 5.688237e-06, 5.728559e-06, 5.721286e-06, 5.733616e-06, 
    5.745416e-06, 5.765227e-06, 5.761967e-06, 5.770697e-06, 5.733298e-06, 
    5.758143e-06, 5.717143e-06, 5.728347e-06, 5.639349e-06, 5.605597e-06, 
    5.591234e-06, 5.578701e-06, 5.548213e-06, 5.56926e-06, 5.56096e-06, 
    5.580721e-06, 5.593283e-06, 5.587071e-06, 5.625457e-06, 5.610523e-06, 
    5.689304e-06, 5.655333e-06, 5.744039e-06, 5.72278e-06, 5.749139e-06, 
    5.735686e-06, 5.758739e-06, 5.737991e-06, 5.773951e-06, 5.781784e-06, 
    5.77643e-06, 5.797019e-06, 5.73684e-06, 5.759926e-06, 5.586895e-06, 
    5.587908e-06, 5.592632e-06, 5.571875e-06, 5.570608e-06, 5.55162e-06, 
    5.568519e-06, 5.575716e-06, 5.594015e-06, 5.604839e-06, 5.615137e-06, 
    5.637798e-06, 5.66313e-06, 5.698618e-06, 5.724157e-06, 5.741291e-06, 
    5.730786e-06, 5.74006e-06, 5.729691e-06, 5.724835e-06, 5.778846e-06, 
    5.748498e-06, 5.794057e-06, 5.791534e-06, 5.770903e-06, 5.791819e-06, 
    5.58862e-06, 5.582791e-06, 5.562554e-06, 5.578389e-06, 5.549553e-06, 
    5.565684e-06, 5.574962e-06, 5.610827e-06, 5.618725e-06, 5.626038e-06, 
    5.640501e-06, 5.659071e-06, 5.691688e-06, 5.720114e-06, 5.746104e-06, 
    5.744199e-06, 5.74487e-06, 5.750675e-06, 5.736292e-06, 5.753038e-06, 
    5.755846e-06, 5.748499e-06, 5.791196e-06, 5.77899e-06, 5.791481e-06, 
    5.783533e-06, 5.584686e-06, 5.594498e-06, 5.589195e-06, 5.599166e-06, 
    5.592138e-06, 5.623398e-06, 5.63278e-06, 5.67675e-06, 5.658703e-06, 
    5.687445e-06, 5.661624e-06, 5.666194e-06, 5.688365e-06, 5.663021e-06, 
    5.718538e-06, 5.680869e-06, 5.750901e-06, 5.71321e-06, 5.753264e-06, 
    5.745992e-06, 5.758038e-06, 5.768829e-06, 5.782419e-06, 5.807505e-06, 
    5.801695e-06, 5.822698e-06, 5.609138e-06, 5.621877e-06, 5.620763e-06, 
    5.634108e-06, 5.643982e-06, 5.665408e-06, 5.699812e-06, 5.686871e-06, 
    5.710644e-06, 5.715417e-06, 5.679307e-06, 5.701463e-06, 5.630414e-06, 
    5.641868e-06, 5.635053e-06, 5.610138e-06, 5.689842e-06, 5.648893e-06, 
    5.724577e-06, 5.702349e-06, 5.767289e-06, 5.734961e-06, 5.798496e-06, 
    5.825693e-06, 5.851356e-06, 5.881341e-06, 5.628842e-06, 5.620181e-06, 
    5.635698e-06, 5.657173e-06, 5.677141e-06, 5.703703e-06, 5.706427e-06, 
    5.711406e-06, 5.724316e-06, 5.735174e-06, 5.712973e-06, 5.737897e-06, 
    5.644511e-06, 5.693404e-06, 5.616901e-06, 5.639896e-06, 5.655909e-06, 
    5.648891e-06, 5.685395e-06, 5.694004e-06, 5.729026e-06, 5.710919e-06, 
    5.81897e-06, 5.771098e-06, 5.904225e-06, 5.866937e-06, 5.617154e-06, 
    5.628815e-06, 5.669444e-06, 5.650104e-06, 5.705482e-06, 5.719132e-06, 
    5.730242e-06, 5.744439e-06, 5.745978e-06, 5.754397e-06, 5.740603e-06, 
    5.753855e-06, 5.70376e-06, 5.726132e-06, 5.664805e-06, 5.679711e-06, 
    5.672855e-06, 5.665332e-06, 5.688559e-06, 5.71332e-06, 5.713862e-06, 
    5.721805e-06, 5.744185e-06, 5.705707e-06, 5.825133e-06, 5.751279e-06, 
    5.641539e-06, 5.664018e-06, 5.667245e-06, 5.658531e-06, 5.717763e-06, 
    5.69628e-06, 5.754193e-06, 5.738528e-06, 5.764204e-06, 5.75144e-06, 
    5.749562e-06, 5.733185e-06, 5.722991e-06, 5.697262e-06, 5.676354e-06, 
    5.659796e-06, 5.663646e-06, 5.68184e-06, 5.714839e-06, 5.746112e-06, 
    5.739256e-06, 5.762251e-06, 5.701461e-06, 5.726924e-06, 5.717075e-06, 
    5.742768e-06, 5.686525e-06, 5.734372e-06, 5.674307e-06, 5.679569e-06, 
    5.695854e-06, 5.728644e-06, 5.735924e-06, 5.743677e-06, 5.738895e-06, 
    5.715679e-06, 5.711883e-06, 5.695461e-06, 5.690923e-06, 5.678425e-06, 
    5.668076e-06, 5.677528e-06, 5.687455e-06, 5.715694e-06, 5.741168e-06, 
    5.76898e-06, 5.775797e-06, 5.808318e-06, 5.781824e-06, 5.825543e-06, 
    5.788343e-06, 5.852792e-06, 5.737167e-06, 5.787274e-06, 5.6966e-06, 
    5.706352e-06, 5.723991e-06, 5.764529e-06, 5.742647e-06, 5.768246e-06, 
    5.711736e-06, 5.682462e-06, 5.674908e-06, 5.6608e-06, 5.675231e-06, 
    5.674057e-06, 5.687875e-06, 5.683435e-06, 5.716632e-06, 5.698794e-06, 
    5.749512e-06, 5.768047e-06, 5.820491e-06, 5.852695e-06, 5.885543e-06, 
    5.900053e-06, 5.904472e-06, 5.906319e-06,
  6.000897e-06, 6.03294e-06, 6.026709e-06, 6.052581e-06, 6.038228e-06, 
    6.055173e-06, 6.007393e-06, 6.03421e-06, 6.017088e-06, 6.003785e-06, 
    6.102883e-06, 6.053738e-06, 6.154107e-06, 6.122657e-06, 6.20177e-06, 
    6.149205e-06, 6.212388e-06, 6.200261e-06, 6.236806e-06, 6.22633e-06, 
    6.273128e-06, 6.241643e-06, 6.297445e-06, 6.26561e-06, 6.270583e-06, 
    6.240604e-06, 6.063626e-06, 6.096755e-06, 6.061663e-06, 6.066383e-06, 
    6.064267e-06, 6.038521e-06, 6.025555e-06, 5.998456e-06, 6.003374e-06, 
    6.023282e-06, 6.068507e-06, 6.053148e-06, 6.091896e-06, 6.091021e-06, 
    6.134245e-06, 6.114744e-06, 6.187548e-06, 6.166831e-06, 6.226768e-06, 
    6.211676e-06, 6.226057e-06, 6.221696e-06, 6.226114e-06, 6.203985e-06, 
    6.213462e-06, 6.194004e-06, 6.118393e-06, 6.140581e-06, 6.074478e-06, 
    6.034832e-06, 6.008566e-06, 5.989945e-06, 5.992576e-06, 5.997592e-06, 
    6.023399e-06, 6.047704e-06, 6.066245e-06, 6.078656e-06, 6.090895e-06, 
    6.127965e-06, 6.147636e-06, 6.191736e-06, 6.183778e-06, 6.197268e-06, 
    6.210175e-06, 6.231854e-06, 6.228285e-06, 6.23784e-06, 6.196918e-06, 
    6.224102e-06, 6.179244e-06, 6.191502e-06, 6.094193e-06, 6.057292e-06, 
    6.041604e-06, 6.027905e-06, 5.994599e-06, 6.017591e-06, 6.008524e-06, 
    6.03011e-06, 6.043836e-06, 6.037048e-06, 6.078996e-06, 6.062675e-06, 
    6.148802e-06, 6.111656e-06, 6.208669e-06, 6.185412e-06, 6.214249e-06, 
    6.19953e-06, 6.224754e-06, 6.202052e-06, 6.2414e-06, 6.249975e-06, 
    6.244114e-06, 6.266648e-06, 6.200793e-06, 6.226054e-06, 6.036856e-06, 
    6.037963e-06, 6.043123e-06, 6.020449e-06, 6.019064e-06, 5.99832e-06, 
    6.016779e-06, 6.024644e-06, 6.044635e-06, 6.056464e-06, 6.067718e-06, 
    6.092486e-06, 6.120182e-06, 6.158986e-06, 6.186918e-06, 6.205662e-06, 
    6.194168e-06, 6.204315e-06, 6.192971e-06, 6.187658e-06, 6.246759e-06, 
    6.213549e-06, 6.263405e-06, 6.260644e-06, 6.238066e-06, 6.260955e-06, 
    6.038741e-06, 6.032371e-06, 6.010264e-06, 6.027562e-06, 5.996063e-06, 
    6.013684e-06, 6.023823e-06, 6.063009e-06, 6.071638e-06, 6.079632e-06, 
    6.095439e-06, 6.115741e-06, 6.151407e-06, 6.182497e-06, 6.210927e-06, 
    6.208843e-06, 6.209577e-06, 6.21593e-06, 6.200193e-06, 6.218515e-06, 
    6.221589e-06, 6.213549e-06, 6.260274e-06, 6.246914e-06, 6.260585e-06, 
    6.251887e-06, 6.034442e-06, 6.045163e-06, 6.039369e-06, 6.050265e-06, 
    6.042586e-06, 6.07675e-06, 6.087005e-06, 6.135075e-06, 6.11534e-06, 
    6.146767e-06, 6.118532e-06, 6.12353e-06, 6.14778e-06, 6.120059e-06, 
    6.180776e-06, 6.13958e-06, 6.216177e-06, 6.174951e-06, 6.218763e-06, 
    6.210804e-06, 6.223986e-06, 6.235795e-06, 6.250667e-06, 6.27813e-06, 
    6.271769e-06, 6.294761e-06, 6.061161e-06, 6.075086e-06, 6.073865e-06, 
    6.088452e-06, 6.099246e-06, 6.122669e-06, 6.160291e-06, 6.146137e-06, 
    6.172136e-06, 6.177358e-06, 6.137866e-06, 6.162098e-06, 6.084416e-06, 
    6.096939e-06, 6.089485e-06, 6.062256e-06, 6.14939e-06, 6.104618e-06, 
    6.187379e-06, 6.163065e-06, 6.23411e-06, 6.19874e-06, 6.268266e-06, 
    6.298047e-06, 6.326142e-06, 6.358992e-06, 6.082696e-06, 6.073229e-06, 
    6.090189e-06, 6.113669e-06, 6.135498e-06, 6.164546e-06, 6.167524e-06, 
    6.17297e-06, 6.187091e-06, 6.198969e-06, 6.174687e-06, 6.201948e-06, 
    6.099833e-06, 6.153283e-06, 6.069646e-06, 6.094784e-06, 6.112286e-06, 
    6.104613e-06, 6.144522e-06, 6.153938e-06, 6.192246e-06, 6.172437e-06, 
    6.290687e-06, 6.238282e-06, 6.384058e-06, 6.343212e-06, 6.069921e-06, 
    6.082666e-06, 6.127084e-06, 6.105938e-06, 6.16649e-06, 6.181422e-06, 
    6.193573e-06, 6.209108e-06, 6.210791e-06, 6.220002e-06, 6.204909e-06, 
    6.219408e-06, 6.164608e-06, 6.189079e-06, 6.122008e-06, 6.138309e-06, 
    6.13081e-06, 6.122585e-06, 6.147983e-06, 6.175067e-06, 6.175656e-06, 
    6.184348e-06, 6.208844e-06, 6.166737e-06, 6.297443e-06, 6.216604e-06, 
    6.096574e-06, 6.121154e-06, 6.124678e-06, 6.11515e-06, 6.179924e-06, 
    6.156428e-06, 6.219779e-06, 6.202639e-06, 6.230733e-06, 6.216767e-06, 
    6.214712e-06, 6.196793e-06, 6.185643e-06, 6.157502e-06, 6.134638e-06, 
    6.116532e-06, 6.120742e-06, 6.140637e-06, 6.176728e-06, 6.210938e-06, 
    6.203438e-06, 6.228596e-06, 6.162094e-06, 6.189947e-06, 6.179174e-06, 
    6.207279e-06, 6.145759e-06, 6.198105e-06, 6.132398e-06, 6.138152e-06, 
    6.155962e-06, 6.191831e-06, 6.19979e-06, 6.208274e-06, 6.20304e-06, 
    6.177647e-06, 6.173494e-06, 6.155531e-06, 6.150569e-06, 6.1369e-06, 
    6.125586e-06, 6.135921e-06, 6.146778e-06, 6.177661e-06, 6.20553e-06, 
    6.235961e-06, 6.24342e-06, 6.279026e-06, 6.250024e-06, 6.297892e-06, 
    6.257169e-06, 6.327726e-06, 6.201158e-06, 6.25599e-06, 6.156776e-06, 
    6.167442e-06, 6.18674e-06, 6.231094e-06, 6.207147e-06, 6.235161e-06, 
    6.173331e-06, 6.141319e-06, 6.133056e-06, 6.117631e-06, 6.133409e-06, 
    6.132125e-06, 6.147234e-06, 6.142378e-06, 6.178687e-06, 6.159176e-06, 
    6.214658e-06, 6.234942e-06, 6.292347e-06, 6.327612e-06, 6.363588e-06, 
    6.379486e-06, 6.384328e-06, 6.386352e-06,
  6.364546e-06, 6.399158e-06, 6.392425e-06, 6.420383e-06, 6.40487e-06, 
    6.423184e-06, 6.371559e-06, 6.400532e-06, 6.382031e-06, 6.367661e-06, 
    6.474778e-06, 6.421633e-06, 6.530194e-06, 6.496156e-06, 6.581805e-06, 
    6.524891e-06, 6.593307e-06, 6.580166e-06, 6.619762e-06, 6.608409e-06, 
    6.659151e-06, 6.625005e-06, 6.685523e-06, 6.650993e-06, 6.656388e-06, 
    6.623879e-06, 6.432318e-06, 6.46815e-06, 6.430196e-06, 6.4353e-06, 
    6.43301e-06, 6.405188e-06, 6.391183e-06, 6.361907e-06, 6.367218e-06, 
    6.388725e-06, 6.437596e-06, 6.420993e-06, 6.462881e-06, 6.461934e-06, 
    6.508694e-06, 6.487594e-06, 6.566397e-06, 6.543961e-06, 6.608882e-06, 
    6.592531e-06, 6.608113e-06, 6.603388e-06, 6.608175e-06, 6.5842e-06, 
    6.594467e-06, 6.573388e-06, 6.491542e-06, 6.515551e-06, 6.444051e-06, 
    6.401208e-06, 6.372828e-06, 6.352717e-06, 6.355558e-06, 6.360975e-06, 
    6.388851e-06, 6.415108e-06, 6.435147e-06, 6.448565e-06, 6.461798e-06, 
    6.501908e-06, 6.52319e-06, 6.570935e-06, 6.562312e-06, 6.576925e-06, 
    6.590905e-06, 6.614396e-06, 6.610528e-06, 6.620885e-06, 6.576543e-06, 
    6.605998e-06, 6.557401e-06, 6.570678e-06, 6.465381e-06, 6.425471e-06, 
    6.408524e-06, 6.393718e-06, 6.357743e-06, 6.382576e-06, 6.372782e-06, 
    6.396097e-06, 6.410929e-06, 6.403593e-06, 6.448932e-06, 6.431289e-06, 
    6.524452e-06, 6.484256e-06, 6.589273e-06, 6.564082e-06, 6.595318e-06, 
    6.579372e-06, 6.606703e-06, 6.582104e-06, 6.624743e-06, 6.63404e-06, 
    6.627686e-06, 6.652114e-06, 6.580741e-06, 6.608112e-06, 6.403387e-06, 
    6.404583e-06, 6.410158e-06, 6.385663e-06, 6.384167e-06, 6.36176e-06, 
    6.381697e-06, 6.390194e-06, 6.41179e-06, 6.424576e-06, 6.43674e-06, 
    6.46352e-06, 6.49348e-06, 6.535473e-06, 6.565714e-06, 6.586014e-06, 
    6.573564e-06, 6.584556e-06, 6.572268e-06, 6.566514e-06, 6.630555e-06, 
    6.594562e-06, 6.648599e-06, 6.645605e-06, 6.621131e-06, 6.645942e-06, 
    6.405422e-06, 6.39854e-06, 6.374661e-06, 6.393345e-06, 6.359322e-06, 
    6.378355e-06, 6.389309e-06, 6.431654e-06, 6.440977e-06, 6.449622e-06, 
    6.466713e-06, 6.488673e-06, 6.527269e-06, 6.560927e-06, 6.591719e-06, 
    6.589461e-06, 6.590256e-06, 6.59714e-06, 6.580091e-06, 6.599941e-06, 
    6.603274e-06, 6.59456e-06, 6.645203e-06, 6.630719e-06, 6.645541e-06, 
    6.636109e-06, 6.400777e-06, 6.412363e-06, 6.406101e-06, 6.417878e-06, 
    6.409579e-06, 6.446509e-06, 6.457599e-06, 6.509596e-06, 6.48824e-06, 
    6.522247e-06, 6.491692e-06, 6.4971e-06, 6.523351e-06, 6.493342e-06, 
    6.559067e-06, 6.514473e-06, 6.597407e-06, 6.552764e-06, 6.600209e-06, 
    6.591586e-06, 6.605868e-06, 6.618668e-06, 6.634788e-06, 6.66457e-06, 
    6.657669e-06, 6.682609e-06, 6.429653e-06, 6.444708e-06, 6.443385e-06, 
    6.459157e-06, 6.470831e-06, 6.496166e-06, 6.536884e-06, 6.521561e-06, 
    6.549705e-06, 6.55536e-06, 6.512609e-06, 6.538841e-06, 6.454795e-06, 
    6.46834e-06, 6.460276e-06, 6.430839e-06, 6.525087e-06, 6.476646e-06, 
    6.566213e-06, 6.539886e-06, 6.616841e-06, 6.578522e-06, 6.653871e-06, 
    6.686181e-06, 6.716662e-06, 6.752337e-06, 6.452934e-06, 6.442697e-06, 
    6.461035e-06, 6.486435e-06, 6.510049e-06, 6.54149e-06, 6.544712e-06, 
    6.55061e-06, 6.565899e-06, 6.578764e-06, 6.552472e-06, 6.581991e-06, 
    6.471478e-06, 6.529299e-06, 6.438826e-06, 6.466011e-06, 6.484938e-06, 
    6.476635e-06, 6.519812e-06, 6.530004e-06, 6.571487e-06, 6.550031e-06, 
    6.678198e-06, 6.621369e-06, 6.77956e-06, 6.735199e-06, 6.439121e-06, 
    6.4529e-06, 6.500947e-06, 6.478069e-06, 6.543593e-06, 6.559761e-06, 
    6.57292e-06, 6.589751e-06, 6.591571e-06, 6.601553e-06, 6.585199e-06, 
    6.600908e-06, 6.541557e-06, 6.568053e-06, 6.495452e-06, 6.51309e-06, 
    6.504974e-06, 6.496075e-06, 6.523558e-06, 6.552885e-06, 6.553517e-06, 
    6.562932e-06, 6.589482e-06, 6.543859e-06, 6.685538e-06, 6.597888e-06, 
    6.46794e-06, 6.494533e-06, 6.498341e-06, 6.488031e-06, 6.558139e-06, 
    6.532701e-06, 6.60131e-06, 6.58274e-06, 6.61318e-06, 6.598046e-06, 
    6.595821e-06, 6.576408e-06, 6.564332e-06, 6.533865e-06, 6.509119e-06, 
    6.489527e-06, 6.49408e-06, 6.515611e-06, 6.554682e-06, 6.591733e-06, 
    6.58361e-06, 6.610864e-06, 6.538833e-06, 6.568996e-06, 6.55733e-06, 
    6.587767e-06, 6.521154e-06, 6.577846e-06, 6.506692e-06, 6.512919e-06, 
    6.532196e-06, 6.57104e-06, 6.579654e-06, 6.588847e-06, 6.583175e-06, 
    6.555676e-06, 6.551177e-06, 6.531729e-06, 6.526361e-06, 6.511564e-06, 
    6.499321e-06, 6.510506e-06, 6.522258e-06, 6.555689e-06, 6.585874e-06, 
    6.618849e-06, 6.626932e-06, 6.665551e-06, 6.6341e-06, 6.686027e-06, 
    6.64186e-06, 6.718396e-06, 6.581146e-06, 6.640571e-06, 6.533076e-06, 
    6.544623e-06, 6.565526e-06, 6.613579e-06, 6.587624e-06, 6.617985e-06, 
    6.551001e-06, 6.516352e-06, 6.507405e-06, 6.490716e-06, 6.507786e-06, 
    6.506397e-06, 6.522748e-06, 6.517492e-06, 6.5568e-06, 6.535674e-06, 
    6.595764e-06, 6.617746e-06, 6.679992e-06, 6.718264e-06, 6.757321e-06, 
    6.77459e-06, 6.779851e-06, 6.78205e-06,
  6.298019e-06, 6.333518e-06, 6.326609e-06, 6.355305e-06, 6.339378e-06, 
    6.358181e-06, 6.305208e-06, 6.33493e-06, 6.315946e-06, 6.30121e-06, 
    6.411204e-06, 6.356588e-06, 6.468217e-06, 6.433178e-06, 6.521402e-06, 
    6.462758e-06, 6.533264e-06, 6.519707e-06, 6.56056e-06, 6.548841e-06, 
    6.601255e-06, 6.565973e-06, 6.628519e-06, 6.592819e-06, 6.598396e-06, 
    6.564811e-06, 6.367557e-06, 6.40439e-06, 6.365379e-06, 6.370623e-06, 
    6.368269e-06, 6.339706e-06, 6.32534e-06, 6.29531e-06, 6.300756e-06, 
    6.322814e-06, 6.372982e-06, 6.355927e-06, 6.398958e-06, 6.397984e-06, 
    6.446079e-06, 6.424369e-06, 6.505511e-06, 6.48239e-06, 6.54933e-06, 
    6.532459e-06, 6.548537e-06, 6.543659e-06, 6.548601e-06, 6.523867e-06, 
    6.534457e-06, 6.512717e-06, 6.428431e-06, 6.453138e-06, 6.37961e-06, 
    6.335629e-06, 6.306509e-06, 6.285892e-06, 6.288804e-06, 6.294358e-06, 
    6.322944e-06, 6.349886e-06, 6.370462e-06, 6.384246e-06, 6.397845e-06, 
    6.439105e-06, 6.461005e-06, 6.510191e-06, 6.5013e-06, 6.516368e-06, 
    6.530782e-06, 6.555022e-06, 6.551029e-06, 6.561721e-06, 6.51597e-06, 
    6.546356e-06, 6.496237e-06, 6.509923e-06, 6.401544e-06, 6.360526e-06, 
    6.343136e-06, 6.327937e-06, 6.291044e-06, 6.316508e-06, 6.306463e-06, 
    6.330376e-06, 6.345597e-06, 6.338066e-06, 6.384623e-06, 6.3665e-06, 
    6.462303e-06, 6.420939e-06, 6.529099e-06, 6.503124e-06, 6.535334e-06, 
    6.518887e-06, 6.547083e-06, 6.521704e-06, 6.565703e-06, 6.575307e-06, 
    6.568743e-06, 6.593975e-06, 6.520298e-06, 6.548537e-06, 6.337855e-06, 
    6.339083e-06, 6.344805e-06, 6.319674e-06, 6.318139e-06, 6.295161e-06, 
    6.315604e-06, 6.324321e-06, 6.346479e-06, 6.359607e-06, 6.3721e-06, 
    6.399616e-06, 6.430427e-06, 6.473651e-06, 6.504806e-06, 6.525737e-06, 
    6.512898e-06, 6.524232e-06, 6.511562e-06, 6.505629e-06, 6.571707e-06, 
    6.534557e-06, 6.590343e-06, 6.587249e-06, 6.561976e-06, 6.587597e-06, 
    6.339945e-06, 6.332881e-06, 6.308388e-06, 6.327551e-06, 6.292662e-06, 
    6.312178e-06, 6.323416e-06, 6.366879e-06, 6.376451e-06, 6.385334e-06, 
    6.402898e-06, 6.425479e-06, 6.465201e-06, 6.499875e-06, 6.53162e-06, 
    6.529292e-06, 6.530111e-06, 6.537214e-06, 6.519629e-06, 6.540104e-06, 
    6.543544e-06, 6.534552e-06, 6.586835e-06, 6.571874e-06, 6.587183e-06, 
    6.57744e-06, 6.335177e-06, 6.347068e-06, 6.340641e-06, 6.35273e-06, 
    6.344212e-06, 6.382139e-06, 6.393535e-06, 6.447011e-06, 6.425034e-06, 
    6.460032e-06, 6.428584e-06, 6.43415e-06, 6.461176e-06, 6.430281e-06, 
    6.49796e-06, 6.452033e-06, 6.53749e-06, 6.491469e-06, 6.540381e-06, 
    6.531483e-06, 6.546219e-06, 6.559432e-06, 6.576076e-06, 6.606851e-06, 
    6.599718e-06, 6.625502e-06, 6.364819e-06, 6.380287e-06, 6.378924e-06, 
    6.395131e-06, 6.407132e-06, 6.433187e-06, 6.475101e-06, 6.459322e-06, 
    6.488307e-06, 6.494135e-06, 6.450106e-06, 6.477119e-06, 6.39065e-06, 
    6.404576e-06, 6.396282e-06, 6.36604e-06, 6.462956e-06, 6.413115e-06, 
    6.505321e-06, 6.478193e-06, 6.557547e-06, 6.518015e-06, 6.595793e-06, 
    6.629204e-06, 6.660737e-06, 6.697698e-06, 6.388737e-06, 6.378217e-06, 
    6.39706e-06, 6.423182e-06, 6.447473e-06, 6.479846e-06, 6.483163e-06, 
    6.489241e-06, 6.504996e-06, 6.51826e-06, 6.491163e-06, 6.521588e-06, 
    6.407809e-06, 6.467292e-06, 6.374243e-06, 6.402182e-06, 6.42164e-06, 
    6.4131e-06, 6.45752e-06, 6.468014e-06, 6.510759e-06, 6.488643e-06, 
    6.620949e-06, 6.562225e-06, 6.725919e-06, 6.67994e-06, 6.374544e-06, 
    6.388701e-06, 6.438109e-06, 6.414574e-06, 6.48201e-06, 6.498671e-06, 
    6.512233e-06, 6.529593e-06, 6.531469e-06, 6.541768e-06, 6.524896e-06, 
    6.541101e-06, 6.479915e-06, 6.507217e-06, 6.43245e-06, 6.450603e-06, 
    6.442248e-06, 6.433092e-06, 6.461377e-06, 6.491588e-06, 6.492235e-06, 
    6.50194e-06, 6.529333e-06, 6.482285e-06, 6.62855e-06, 6.538002e-06, 
    6.404158e-06, 6.431513e-06, 6.435425e-06, 6.424817e-06, 6.497e-06, 
    6.470793e-06, 6.541517e-06, 6.52236e-06, 6.553765e-06, 6.538149e-06, 
    6.535853e-06, 6.51583e-06, 6.503382e-06, 6.471993e-06, 6.446517e-06, 
    6.426355e-06, 6.43104e-06, 6.453199e-06, 6.49344e-06, 6.531639e-06, 
    6.52326e-06, 6.551375e-06, 6.477108e-06, 6.508191e-06, 6.496168e-06, 
    6.527545e-06, 6.458903e-06, 6.51733e-06, 6.444016e-06, 6.450426e-06, 
    6.470274e-06, 6.510302e-06, 6.519177e-06, 6.528661e-06, 6.522808e-06, 
    6.494463e-06, 6.489825e-06, 6.469791e-06, 6.464265e-06, 6.44903e-06, 
    6.436432e-06, 6.447941e-06, 6.460042e-06, 6.494474e-06, 6.525595e-06, 
    6.55962e-06, 6.567962e-06, 6.607875e-06, 6.575375e-06, 6.629057e-06, 
    6.583402e-06, 6.662548e-06, 6.520725e-06, 6.58206e-06, 6.471177e-06, 
    6.483071e-06, 6.504617e-06, 6.554184e-06, 6.527398e-06, 6.558731e-06, 
    6.489644e-06, 6.453964e-06, 6.44475e-06, 6.427581e-06, 6.445143e-06, 
    6.443714e-06, 6.460542e-06, 6.455132e-06, 6.49562e-06, 6.473854e-06, 
    6.535795e-06, 6.558483e-06, 6.622797e-06, 6.662402e-06, 6.702856e-06, 
    6.720762e-06, 6.726217e-06, 6.728499e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.777233, 5.777218, 5.777221, 5.777209, 5.777215, 5.777208, 5.77723, 
    5.777217, 5.777225, 5.777231, 5.777186, 5.777208, 5.777163, 5.777177, 
    5.777142, 5.777165, 5.777137, 5.777142, 5.777126, 5.77713, 5.777109, 
    5.777123, 5.777098, 5.777112, 5.777111, 5.777124, 5.777204, 5.777189, 
    5.777205, 5.777203, 5.777204, 5.777215, 5.777221, 5.777234, 5.777231, 
    5.777222, 5.777202, 5.777209, 5.777191, 5.777192, 5.777172, 5.777181, 
    5.777148, 5.777157, 5.77713, 5.777137, 5.777131, 5.777133, 5.777131, 
    5.777141, 5.777136, 5.777145, 5.777179, 5.777169, 5.777199, 5.777217, 
    5.777229, 5.777237, 5.777236, 5.777234, 5.777222, 5.777211, 5.777203, 
    5.777197, 5.777192, 5.777175, 5.777166, 5.777146, 5.77715, 5.777143, 
    5.777138, 5.777128, 5.77713, 5.777125, 5.777143, 5.777132, 5.777152, 
    5.777146, 5.77719, 5.777207, 5.777214, 5.77722, 5.777236, 5.777225, 
    5.777229, 5.777219, 5.777213, 5.777216, 5.777197, 5.777205, 5.777165, 
    5.777182, 5.777138, 5.777149, 5.777136, 5.777143, 5.777131, 5.777141, 
    5.777123, 5.77712, 5.777122, 5.777112, 5.777142, 5.777131, 5.777216, 
    5.777215, 5.777213, 5.777224, 5.777224, 5.777234, 5.777225, 5.777222, 
    5.777213, 5.777207, 5.777202, 5.777191, 5.777178, 5.777161, 5.777148, 
    5.77714, 5.777145, 5.77714, 5.777145, 5.777148, 5.777121, 5.777136, 
    5.777113, 5.777115, 5.777125, 5.777115, 5.777215, 5.777218, 5.777228, 
    5.77722, 5.777235, 5.777227, 5.777222, 5.777204, 5.7772, 5.777197, 
    5.77719, 5.77718, 5.777164, 5.77715, 5.777137, 5.777138, 5.777138, 
    5.777135, 5.777142, 5.777134, 5.777133, 5.777136, 5.777115, 5.777121, 
    5.777115, 5.777119, 5.777217, 5.777212, 5.777215, 5.77721, 5.777214, 
    5.777198, 5.777194, 5.777172, 5.777181, 5.777166, 5.777179, 5.777177, 
    5.777166, 5.777178, 5.777151, 5.77717, 5.777135, 5.777153, 5.777134, 
    5.777137, 5.777132, 5.777126, 5.777119, 5.777107, 5.77711, 5.7771, 
    5.777205, 5.777199, 5.777199, 5.777193, 5.777188, 5.777177, 5.77716, 
    5.777166, 5.777155, 5.777153, 5.77717, 5.777159, 5.777194, 5.777189, 
    5.777192, 5.777205, 5.777165, 5.777185, 5.777148, 5.777159, 5.777127, 
    5.777143, 5.777112, 5.777098, 5.777085, 5.777071, 5.777195, 5.7772, 
    5.777192, 5.777181, 5.777171, 5.777158, 5.777157, 5.777154, 5.777148, 
    5.777143, 5.777153, 5.777141, 5.777187, 5.777164, 5.777201, 5.77719, 
    5.777182, 5.777185, 5.777167, 5.777163, 5.777146, 5.777154, 5.777102, 
    5.777125, 5.77706, 5.777078, 5.777201, 5.777195, 5.777175, 5.777185, 
    5.777157, 5.777151, 5.777145, 5.777138, 5.777137, 5.777133, 5.77714, 
    5.777133, 5.777158, 5.777147, 5.777177, 5.77717, 5.777174, 5.777177, 
    5.777166, 5.777153, 5.777153, 5.777149, 5.777138, 5.777157, 5.777098, 
    5.777135, 5.777189, 5.777178, 5.777176, 5.777181, 5.777151, 5.777162, 
    5.777133, 5.777141, 5.777128, 5.777134, 5.777135, 5.777143, 5.777149, 
    5.777162, 5.777172, 5.77718, 5.777178, 5.777169, 5.777153, 5.777137, 
    5.777141, 5.777129, 5.777159, 5.777147, 5.777152, 5.777139, 5.777167, 
    5.777143, 5.777173, 5.77717, 5.777162, 5.777146, 5.777142, 5.777138, 
    5.777141, 5.777152, 5.777154, 5.777162, 5.777164, 5.777171, 5.777176, 
    5.777171, 5.777166, 5.777152, 5.77714, 5.777126, 5.777122, 5.777107, 
    5.77712, 5.777098, 5.777116, 5.777085, 5.777142, 5.777117, 5.777162, 
    5.777157, 5.777148, 5.777128, 5.777139, 5.777126, 5.777154, 5.777169, 
    5.777173, 5.777179, 5.777172, 5.777173, 5.777166, 5.777168, 5.777152, 
    5.777161, 5.777135, 5.777126, 5.777101, 5.777085, 5.777069, 5.777061, 
    5.77706, 5.777059 ;

 SOIL1C_TO_SOIL2C =
  3.814359e-08, 3.824792e-08, 3.822764e-08, 3.831176e-08, 3.826511e-08, 
    3.832018e-08, 3.816475e-08, 3.825205e-08, 3.819632e-08, 3.815299e-08, 
    3.847494e-08, 3.831552e-08, 3.864054e-08, 3.853891e-08, 3.879418e-08, 
    3.862472e-08, 3.882835e-08, 3.878932e-08, 3.890683e-08, 3.887317e-08, 
    3.90234e-08, 3.892237e-08, 3.910128e-08, 3.899929e-08, 3.901523e-08, 
    3.891903e-08, 3.834762e-08, 3.845509e-08, 3.834125e-08, 3.835658e-08, 
    3.83497e-08, 3.826606e-08, 3.82239e-08, 3.813562e-08, 3.815165e-08, 
    3.821649e-08, 3.836347e-08, 3.831359e-08, 3.843931e-08, 3.843648e-08, 
    3.857637e-08, 3.85133e-08, 3.874838e-08, 3.868158e-08, 3.887457e-08, 
    3.882604e-08, 3.887229e-08, 3.885827e-08, 3.887248e-08, 3.88013e-08, 
    3.88318e-08, 3.876917e-08, 3.852511e-08, 3.859685e-08, 3.838284e-08, 
    3.825408e-08, 3.816857e-08, 3.810787e-08, 3.811645e-08, 3.813281e-08, 
    3.821687e-08, 3.829591e-08, 3.835612e-08, 3.839639e-08, 3.843607e-08, 
    3.855609e-08, 3.861965e-08, 3.876187e-08, 3.873622e-08, 3.877968e-08, 
    3.882122e-08, 3.889092e-08, 3.887945e-08, 3.891016e-08, 3.877855e-08, 
    3.886601e-08, 3.872161e-08, 3.876111e-08, 3.84468e-08, 3.832706e-08, 
    3.82761e-08, 3.823153e-08, 3.812305e-08, 3.819797e-08, 3.816843e-08, 
    3.82387e-08, 3.828334e-08, 3.826127e-08, 3.839749e-08, 3.834453e-08, 
    3.862341e-08, 3.850332e-08, 3.881637e-08, 3.874149e-08, 3.883432e-08, 
    3.878696e-08, 3.886811e-08, 3.879508e-08, 3.892159e-08, 3.894912e-08, 
    3.893031e-08, 3.90026e-08, 3.879103e-08, 3.887229e-08, 3.826064e-08, 
    3.826424e-08, 3.828102e-08, 3.820727e-08, 3.820276e-08, 3.813518e-08, 
    3.819532e-08, 3.822092e-08, 3.828593e-08, 3.832437e-08, 3.83609e-08, 
    3.844123e-08, 3.85309e-08, 3.865628e-08, 3.874634e-08, 3.880669e-08, 
    3.876969e-08, 3.880236e-08, 3.876584e-08, 3.874872e-08, 3.89388e-08, 
    3.883208e-08, 3.899221e-08, 3.898335e-08, 3.891088e-08, 3.898435e-08, 
    3.826677e-08, 3.824605e-08, 3.81741e-08, 3.823041e-08, 3.812782e-08, 
    3.818524e-08, 3.821825e-08, 3.834563e-08, 3.837362e-08, 3.839956e-08, 
    3.845079e-08, 3.851653e-08, 3.863182e-08, 3.87321e-08, 3.882364e-08, 
    3.881693e-08, 3.881929e-08, 3.883973e-08, 3.878909e-08, 3.884804e-08, 
    3.885793e-08, 3.883207e-08, 3.898216e-08, 3.893929e-08, 3.898316e-08, 
    3.895525e-08, 3.825279e-08, 3.828765e-08, 3.826881e-08, 3.830423e-08, 
    3.827927e-08, 3.839022e-08, 3.842348e-08, 3.857906e-08, 3.851523e-08, 
    3.861683e-08, 3.852556e-08, 3.854173e-08, 3.862013e-08, 3.853049e-08, 
    3.872656e-08, 3.859363e-08, 3.884053e-08, 3.87078e-08, 3.884884e-08, 
    3.882324e-08, 3.886563e-08, 3.890359e-08, 3.895134e-08, 3.903942e-08, 
    3.901903e-08, 3.909268e-08, 3.833962e-08, 3.838482e-08, 3.838085e-08, 
    3.842815e-08, 3.846313e-08, 3.853894e-08, 3.866049e-08, 3.861479e-08, 
    3.869869e-08, 3.871553e-08, 3.858807e-08, 3.866632e-08, 3.841507e-08, 
    3.845566e-08, 3.84315e-08, 3.834318e-08, 3.862531e-08, 3.848054e-08, 
    3.874783e-08, 3.866944e-08, 3.889817e-08, 3.878443e-08, 3.90078e-08, 
    3.910322e-08, 3.919305e-08, 3.929794e-08, 3.840949e-08, 3.837878e-08, 
    3.843378e-08, 3.850983e-08, 3.858042e-08, 3.867422e-08, 3.868382e-08, 
    3.870139e-08, 3.87469e-08, 3.878515e-08, 3.870693e-08, 3.879474e-08, 
    3.846506e-08, 3.863787e-08, 3.836717e-08, 3.844869e-08, 3.850536e-08, 
    3.848051e-08, 3.860957e-08, 3.863997e-08, 3.876351e-08, 3.869966e-08, 
    3.907966e-08, 3.891159e-08, 3.937783e-08, 3.924759e-08, 3.836805e-08, 
    3.840939e-08, 3.855322e-08, 3.84848e-08, 3.868048e-08, 3.872863e-08, 
    3.876778e-08, 3.881779e-08, 3.88232e-08, 3.885283e-08, 3.880427e-08, 
    3.885091e-08, 3.867442e-08, 3.87533e-08, 3.85368e-08, 3.85895e-08, 
    3.856526e-08, 3.853867e-08, 3.862075e-08, 3.870816e-08, 3.871004e-08, 
    3.873807e-08, 3.881698e-08, 3.868128e-08, 3.910131e-08, 3.884194e-08, 
    3.845447e-08, 3.853405e-08, 3.854544e-08, 3.851461e-08, 3.87238e-08, 
    3.864802e-08, 3.885211e-08, 3.879697e-08, 3.888731e-08, 3.884242e-08, 
    3.883581e-08, 3.877815e-08, 3.874223e-08, 3.865149e-08, 3.857764e-08, 
    3.851909e-08, 3.85327e-08, 3.859703e-08, 3.871351e-08, 3.882368e-08, 
    3.879955e-08, 3.888045e-08, 3.86663e-08, 3.87561e-08, 3.872139e-08, 
    3.88119e-08, 3.861357e-08, 3.878241e-08, 3.857039e-08, 3.858899e-08, 
    3.864652e-08, 3.876218e-08, 3.878779e-08, 3.881511e-08, 3.879826e-08, 
    3.871647e-08, 3.870307e-08, 3.864512e-08, 3.862911e-08, 3.858495e-08, 
    3.854837e-08, 3.858178e-08, 3.861687e-08, 3.871651e-08, 3.880627e-08, 
    3.890412e-08, 3.892807e-08, 3.904231e-08, 3.89493e-08, 3.910275e-08, 
    3.897226e-08, 3.919815e-08, 3.879222e-08, 3.896845e-08, 3.864914e-08, 
    3.868355e-08, 3.874578e-08, 3.888849e-08, 3.881147e-08, 3.890156e-08, 
    3.870255e-08, 3.859924e-08, 3.857252e-08, 3.852264e-08, 3.857366e-08, 
    3.856951e-08, 3.861833e-08, 3.860265e-08, 3.871982e-08, 3.865689e-08, 
    3.883564e-08, 3.890085e-08, 3.908496e-08, 3.919777e-08, 3.931259e-08, 
    3.936326e-08, 3.937868e-08, 3.938513e-08 ;

 SOIL1C_TO_SOIL3C =
  4.523483e-10, 4.535861e-10, 4.533456e-10, 4.543436e-10, 4.537901e-10, 
    4.544435e-10, 4.525994e-10, 4.536352e-10, 4.52974e-10, 4.524599e-10, 
    4.562797e-10, 4.543882e-10, 4.582446e-10, 4.570387e-10, 4.600676e-10, 
    4.580569e-10, 4.60473e-10, 4.600098e-10, 4.614042e-10, 4.610048e-10, 
    4.627873e-10, 4.615885e-10, 4.637114e-10, 4.625012e-10, 4.626904e-10, 
    4.615489e-10, 4.547691e-10, 4.560442e-10, 4.546935e-10, 4.548754e-10, 
    4.547938e-10, 4.538015e-10, 4.533011e-10, 4.522538e-10, 4.52444e-10, 
    4.532133e-10, 4.549572e-10, 4.543654e-10, 4.55857e-10, 4.558234e-10, 
    4.574832e-10, 4.567349e-10, 4.595241e-10, 4.587316e-10, 4.610214e-10, 
    4.604457e-10, 4.609944e-10, 4.60828e-10, 4.609965e-10, 4.601521e-10, 
    4.605138e-10, 4.597707e-10, 4.56875e-10, 4.577262e-10, 4.55187e-10, 
    4.536593e-10, 4.526448e-10, 4.519246e-10, 4.520264e-10, 4.522205e-10, 
    4.532178e-10, 4.541555e-10, 4.548699e-10, 4.553477e-10, 4.558185e-10, 
    4.572426e-10, 4.579967e-10, 4.596842e-10, 4.593799e-10, 4.598955e-10, 
    4.603884e-10, 4.612154e-10, 4.610793e-10, 4.614436e-10, 4.598821e-10, 
    4.609199e-10, 4.592065e-10, 4.596751e-10, 4.559458e-10, 4.545251e-10, 
    4.539205e-10, 4.533918e-10, 4.521047e-10, 4.529935e-10, 4.526431e-10, 
    4.534768e-10, 4.540064e-10, 4.537445e-10, 4.553608e-10, 4.547325e-10, 
    4.580413e-10, 4.566164e-10, 4.603309e-10, 4.594423e-10, 4.605439e-10, 
    4.599819e-10, 4.609447e-10, 4.600782e-10, 4.615793e-10, 4.61906e-10, 
    4.616827e-10, 4.625406e-10, 4.600301e-10, 4.609943e-10, 4.537372e-10, 
    4.537798e-10, 4.539789e-10, 4.531039e-10, 4.530504e-10, 4.522486e-10, 
    4.529621e-10, 4.532658e-10, 4.540371e-10, 4.544932e-10, 4.549267e-10, 
    4.558797e-10, 4.569437e-10, 4.584313e-10, 4.594999e-10, 4.60216e-10, 
    4.59777e-10, 4.601646e-10, 4.597313e-10, 4.595282e-10, 4.617835e-10, 
    4.605172e-10, 4.624172e-10, 4.623121e-10, 4.614523e-10, 4.62324e-10, 
    4.538099e-10, 4.535641e-10, 4.527104e-10, 4.533785e-10, 4.521613e-10, 
    4.528425e-10, 4.532342e-10, 4.547455e-10, 4.550776e-10, 4.553853e-10, 
    4.559932e-10, 4.567732e-10, 4.581411e-10, 4.59331e-10, 4.604171e-10, 
    4.603375e-10, 4.603655e-10, 4.60608e-10, 4.600072e-10, 4.607067e-10, 
    4.60824e-10, 4.605171e-10, 4.62298e-10, 4.617893e-10, 4.623099e-10, 
    4.619787e-10, 4.53644e-10, 4.540576e-10, 4.538341e-10, 4.542543e-10, 
    4.539582e-10, 4.552745e-10, 4.556691e-10, 4.575152e-10, 4.567578e-10, 
    4.579633e-10, 4.568803e-10, 4.570722e-10, 4.580024e-10, 4.569389e-10, 
    4.592652e-10, 4.57688e-10, 4.606174e-10, 4.590426e-10, 4.607161e-10, 
    4.604124e-10, 4.609153e-10, 4.613657e-10, 4.619323e-10, 4.629774e-10, 
    4.627355e-10, 4.636094e-10, 4.546742e-10, 4.552104e-10, 4.551634e-10, 
    4.557246e-10, 4.561396e-10, 4.570391e-10, 4.584813e-10, 4.57939e-10, 
    4.589346e-10, 4.591343e-10, 4.57622e-10, 4.585505e-10, 4.555694e-10, 
    4.56051e-10, 4.557644e-10, 4.547164e-10, 4.580638e-10, 4.563462e-10, 
    4.595176e-10, 4.585875e-10, 4.613014e-10, 4.599518e-10, 4.626022e-10, 
    4.637344e-10, 4.648004e-10, 4.66045e-10, 4.555032e-10, 4.551388e-10, 
    4.557913e-10, 4.566937e-10, 4.575312e-10, 4.586442e-10, 4.587581e-10, 
    4.589665e-10, 4.595065e-10, 4.599604e-10, 4.590323e-10, 4.600742e-10, 
    4.561625e-10, 4.582129e-10, 4.55001e-10, 4.559682e-10, 4.566406e-10, 
    4.563458e-10, 4.578771e-10, 4.582379e-10, 4.597037e-10, 4.589461e-10, 
    4.634549e-10, 4.614606e-10, 4.669929e-10, 4.654475e-10, 4.550115e-10, 
    4.55502e-10, 4.572086e-10, 4.563967e-10, 4.587185e-10, 4.592898e-10, 
    4.597542e-10, 4.603477e-10, 4.604118e-10, 4.607634e-10, 4.601873e-10, 
    4.607407e-10, 4.586465e-10, 4.595825e-10, 4.570137e-10, 4.57639e-10, 
    4.573514e-10, 4.570358e-10, 4.580097e-10, 4.590469e-10, 4.590693e-10, 
    4.594017e-10, 4.603381e-10, 4.587279e-10, 4.637118e-10, 4.606343e-10, 
    4.560368e-10, 4.569811e-10, 4.571162e-10, 4.567504e-10, 4.592325e-10, 
    4.583333e-10, 4.607549e-10, 4.601006e-10, 4.611726e-10, 4.606399e-10, 
    4.605615e-10, 4.598773e-10, 4.594512e-10, 4.583745e-10, 4.574983e-10, 
    4.568035e-10, 4.569651e-10, 4.577283e-10, 4.591104e-10, 4.604175e-10, 
    4.601312e-10, 4.610912e-10, 4.585502e-10, 4.596158e-10, 4.592039e-10, 
    4.602778e-10, 4.579246e-10, 4.599279e-10, 4.574123e-10, 4.57633e-10, 
    4.583155e-10, 4.596879e-10, 4.599918e-10, 4.603158e-10, 4.601159e-10, 
    4.591455e-10, 4.589865e-10, 4.582989e-10, 4.581089e-10, 4.575849e-10, 
    4.57151e-10, 4.575474e-10, 4.579637e-10, 4.59146e-10, 4.602111e-10, 
    4.61372e-10, 4.616562e-10, 4.630117e-10, 4.619081e-10, 4.637289e-10, 
    4.621805e-10, 4.648609e-10, 4.600443e-10, 4.621353e-10, 4.583466e-10, 
    4.58755e-10, 4.594933e-10, 4.611866e-10, 4.602727e-10, 4.613416e-10, 
    4.589804e-10, 4.577546e-10, 4.574375e-10, 4.568457e-10, 4.574511e-10, 
    4.574019e-10, 4.579811e-10, 4.57795e-10, 4.591852e-10, 4.584385e-10, 
    4.605595e-10, 4.613332e-10, 4.635178e-10, 4.648563e-10, 4.662188e-10, 
    4.6682e-10, 4.67003e-10, 4.670795e-10 ;

 SOIL1C_vr =
  19.98041, 19.98036, 19.98037, 19.98033, 19.98035, 19.98033, 19.9804, 
    19.98036, 19.98038, 19.98041, 19.98025, 19.98033, 19.98017, 19.98022, 
    19.9801, 19.98018, 19.98008, 19.9801, 19.98004, 19.98006, 19.97999, 
    19.98004, 19.97995, 19.98, 19.97999, 19.98004, 19.98031, 19.98026, 
    19.98031, 19.98031, 19.98031, 19.98035, 19.98037, 19.98041, 19.98041, 
    19.98038, 19.9803, 19.98033, 19.98027, 19.98027, 19.9802, 19.98023, 
    19.98012, 19.98015, 19.98006, 19.98008, 19.98006, 19.98007, 19.98006, 
    19.98009, 19.98008, 19.98011, 19.98023, 19.98019, 19.9803, 19.98036, 
    19.9804, 19.98043, 19.98042, 19.98042, 19.98038, 19.98034, 19.98031, 
    19.98029, 19.98027, 19.98021, 19.98018, 19.98011, 19.98013, 19.9801, 
    19.98008, 19.98005, 19.98006, 19.98004, 19.9801, 19.98006, 19.98013, 
    19.98011, 19.98026, 19.98032, 19.98035, 19.98037, 19.98042, 19.98038, 
    19.9804, 19.98036, 19.98034, 19.98035, 19.98029, 19.98031, 19.98018, 
    19.98024, 19.98009, 19.98012, 19.98008, 19.9801, 19.98006, 19.9801, 
    19.98004, 19.98002, 19.98003, 19.98, 19.9801, 19.98006, 19.98035, 
    19.98035, 19.98034, 19.98038, 19.98038, 19.98041, 19.98038, 19.98037, 
    19.98034, 19.98032, 19.9803, 19.98027, 19.98022, 19.98016, 19.98012, 
    19.98009, 19.98011, 19.98009, 19.98011, 19.98012, 19.98003, 19.98008, 
    19.98, 19.98001, 19.98004, 19.98001, 19.98035, 19.98036, 19.9804, 
    19.98037, 19.98042, 19.98039, 19.98037, 19.98031, 19.9803, 19.98029, 
    19.98026, 19.98023, 19.98018, 19.98013, 19.98008, 19.98009, 19.98009, 
    19.98008, 19.9801, 19.98007, 19.98007, 19.98008, 19.98001, 19.98003, 
    19.98001, 19.98002, 19.98036, 19.98034, 19.98035, 19.98033, 19.98034, 
    19.98029, 19.98028, 19.9802, 19.98023, 19.98018, 19.98023, 19.98022, 
    19.98018, 19.98022, 19.98013, 19.98019, 19.98008, 19.98014, 19.98007, 
    19.98008, 19.98006, 19.98005, 19.98002, 19.97998, 19.97999, 19.97995, 
    19.98032, 19.98029, 19.9803, 19.98027, 19.98026, 19.98022, 19.98016, 
    19.98018, 19.98014, 19.98013, 19.9802, 19.98016, 19.98028, 19.98026, 
    19.98027, 19.98031, 19.98018, 19.98025, 19.98012, 19.98016, 19.98005, 
    19.9801, 19.98, 19.97995, 19.97991, 19.97986, 19.98028, 19.9803, 
    19.98027, 19.98023, 19.9802, 19.98015, 19.98015, 19.98014, 19.98012, 
    19.9801, 19.98014, 19.9801, 19.98026, 19.98017, 19.9803, 19.98026, 
    19.98024, 19.98025, 19.98019, 19.98017, 19.98011, 19.98014, 19.97996, 
    19.98004, 19.97982, 19.97988, 19.9803, 19.98028, 19.98021, 19.98025, 
    19.98015, 19.98013, 19.98011, 19.98009, 19.98008, 19.98007, 19.98009, 
    19.98007, 19.98015, 19.98012, 19.98022, 19.9802, 19.98021, 19.98022, 
    19.98018, 19.98014, 19.98014, 19.98012, 19.98009, 19.98015, 19.97995, 
    19.98007, 19.98026, 19.98022, 19.98022, 19.98023, 19.98013, 19.98017, 
    19.98007, 19.9801, 19.98005, 19.98007, 19.98008, 19.9801, 19.98012, 
    19.98017, 19.9802, 19.98023, 19.98022, 19.98019, 19.98014, 19.98008, 
    19.98009, 19.98006, 19.98016, 19.98012, 19.98013, 19.98009, 19.98018, 
    19.9801, 19.98021, 19.9802, 19.98017, 19.98011, 19.9801, 19.98009, 
    19.98009, 19.98013, 19.98014, 19.98017, 19.98018, 19.9802, 19.98022, 
    19.9802, 19.98018, 19.98013, 19.98009, 19.98005, 19.98003, 19.97998, 
    19.98002, 19.97995, 19.98001, 19.9799, 19.9801, 19.98001, 19.98017, 
    19.98015, 19.98012, 19.98005, 19.98009, 19.98005, 19.98014, 19.98019, 
    19.9802, 19.98023, 19.9802, 19.98021, 19.98018, 19.98019, 19.98013, 
    19.98016, 19.98008, 19.98005, 19.97996, 19.9799, 19.97985, 19.97983, 
    19.97982, 19.97981,
  19.98022, 19.98017, 19.98018, 19.98014, 19.98016, 19.98013, 19.98021, 
    19.98017, 19.9802, 19.98022, 19.98006, 19.98014, 19.97997, 19.98003, 
    19.9799, 19.97998, 19.97988, 19.9799, 19.97984, 19.97986, 19.97978, 
    19.97984, 19.97975, 19.9798, 19.97979, 19.97984, 19.98012, 19.98007, 
    19.98013, 19.98012, 19.98012, 19.98016, 19.98018, 19.98023, 19.98022, 
    19.98019, 19.98011, 19.98014, 19.98008, 19.98008, 19.98001, 19.98004, 
    19.97992, 19.97996, 19.97986, 19.97988, 19.97986, 19.97987, 19.97986, 
    19.97989, 19.97988, 19.97991, 19.98003, 19.98, 19.9801, 19.98017, 
    19.98021, 19.98024, 19.98024, 19.98023, 19.98019, 19.98015, 19.98012, 
    19.9801, 19.98008, 19.98002, 19.97999, 19.97992, 19.97993, 19.97991, 
    19.97989, 19.97985, 19.97986, 19.97984, 19.97991, 19.97986, 19.97993, 
    19.97992, 19.98007, 19.98013, 19.98016, 19.98018, 19.98023, 19.9802, 
    19.98021, 19.98018, 19.98015, 19.98017, 19.9801, 19.98012, 19.97998, 
    19.98004, 19.97989, 19.97993, 19.97988, 19.9799, 19.97986, 19.9799, 
    19.97984, 19.97982, 19.97983, 19.9798, 19.9799, 19.97986, 19.98017, 
    19.98016, 19.98015, 19.98019, 19.98019, 19.98023, 19.9802, 19.98018, 
    19.98015, 19.98013, 19.98011, 19.98007, 19.98003, 19.97997, 19.97992, 
    19.97989, 19.97991, 19.97989, 19.97991, 19.97992, 19.97983, 19.97988, 
    19.9798, 19.9798, 19.97984, 19.9798, 19.98016, 19.98017, 19.98021, 
    19.98018, 19.98023, 19.9802, 19.98019, 19.98012, 19.98011, 19.98009, 
    19.98007, 19.98004, 19.97998, 19.97993, 19.97988, 19.97989, 19.97989, 
    19.97988, 19.9799, 19.97987, 19.97987, 19.97988, 19.9798, 19.97983, 
    19.9798, 19.97982, 19.98017, 19.98015, 19.98016, 19.98014, 19.98016, 
    19.9801, 19.98008, 19.98001, 19.98004, 19.97999, 19.98003, 19.98002, 
    19.97999, 19.98003, 19.97993, 19.98, 19.97988, 19.97994, 19.97987, 
    19.97989, 19.97986, 19.97985, 19.97982, 19.97978, 19.97979, 19.97975, 
    19.98013, 19.9801, 19.9801, 19.98008, 19.98006, 19.98003, 19.97997, 
    19.97999, 19.97995, 19.97994, 19.98, 19.97996, 19.98009, 19.98007, 
    19.98008, 19.98012, 19.97998, 19.98005, 19.97992, 19.97996, 19.97985, 
    19.9799, 19.97979, 19.97975, 19.9797, 19.97965, 19.98009, 19.98011, 
    19.98008, 19.98004, 19.98001, 19.97996, 19.97995, 19.97994, 19.97992, 
    19.9799, 19.97994, 19.9799, 19.98006, 19.97998, 19.98011, 19.98007, 
    19.98004, 19.98005, 19.97999, 19.97997, 19.97991, 19.97995, 19.97976, 
    19.97984, 19.97961, 19.97967, 19.98011, 19.98009, 19.98002, 19.98005, 
    19.97996, 19.97993, 19.97991, 19.97989, 19.97989, 19.97987, 19.97989, 
    19.97987, 19.97996, 19.97992, 19.98003, 19.98, 19.98001, 19.98003, 
    19.97998, 19.97994, 19.97994, 19.97993, 19.97989, 19.97996, 19.97975, 
    19.97988, 19.98007, 19.98003, 19.98002, 19.98004, 19.97993, 19.97997, 
    19.97987, 19.9799, 19.97985, 19.97988, 19.97988, 19.97991, 19.97993, 
    19.97997, 19.98001, 19.98004, 19.98003, 19.98, 19.97994, 19.97988, 
    19.9799, 19.97986, 19.97996, 19.97992, 19.97993, 19.97989, 19.97999, 
    19.9799, 19.98001, 19.98, 19.97997, 19.97991, 19.9799, 19.97989, 19.9799, 
    19.97994, 19.97994, 19.97997, 19.97998, 19.98, 19.98002, 19.98001, 
    19.97999, 19.97994, 19.97989, 19.97984, 19.97983, 19.97977, 19.97982, 
    19.97975, 19.97981, 19.9797, 19.9799, 19.97981, 19.97997, 19.97995, 
    19.97992, 19.97985, 19.97989, 19.97985, 19.97994, 19.98, 19.98001, 
    19.98003, 19.98001, 19.98001, 19.97999, 19.97999, 19.97994, 19.97997, 
    19.97988, 19.97985, 19.97975, 19.9797, 19.97964, 19.97962, 19.97961, 
    19.9796,
  19.98016, 19.98011, 19.98012, 19.98007, 19.9801, 19.98007, 19.98015, 
    19.9801, 19.98013, 19.98015, 19.97999, 19.98007, 19.97991, 19.97996, 
    19.97983, 19.97992, 19.97981, 19.97983, 19.97977, 19.97979, 19.97971, 
    19.97976, 19.97967, 19.97972, 19.97972, 19.97977, 19.98005, 19.98, 
    19.98006, 19.98005, 19.98005, 19.9801, 19.98012, 19.98016, 19.98015, 
    19.98012, 19.98005, 19.98007, 19.98001, 19.98001, 19.97994, 19.97997, 
    19.97985, 19.97989, 19.97979, 19.97981, 19.97979, 19.9798, 19.97979, 
    19.97983, 19.97981, 19.97984, 19.97997, 19.97993, 19.98004, 19.9801, 
    19.98015, 19.98018, 19.98017, 19.98016, 19.98012, 19.98008, 19.98005, 
    19.98003, 19.98001, 19.97995, 19.97992, 19.97985, 19.97986, 19.97984, 
    19.97982, 19.97978, 19.97979, 19.97977, 19.97984, 19.97979, 19.97987, 
    19.97985, 19.98001, 19.98007, 19.98009, 19.98011, 19.98017, 19.98013, 
    19.98015, 19.98011, 19.98009, 19.9801, 19.98003, 19.98006, 19.97992, 
    19.97998, 19.97982, 19.97986, 19.97981, 19.97983, 19.97979, 19.97983, 
    19.97976, 19.97975, 19.97976, 19.97972, 19.97983, 19.97979, 19.9801, 
    19.9801, 19.98009, 19.98013, 19.98013, 19.98016, 19.98013, 19.98012, 
    19.98009, 19.98007, 19.98005, 19.98001, 19.97996, 19.9799, 19.97985, 
    19.97982, 19.97984, 19.97983, 19.97984, 19.97985, 19.97976, 19.97981, 
    19.97973, 19.97973, 19.97977, 19.97973, 19.9801, 19.98011, 19.98014, 
    19.98011, 19.98017, 19.98014, 19.98012, 19.98006, 19.98004, 19.98003, 
    19.98, 19.97997, 19.97991, 19.97986, 19.97981, 19.97982, 19.97982, 
    19.97981, 19.97983, 19.9798, 19.9798, 19.97981, 19.97973, 19.97976, 
    19.97973, 19.97975, 19.9801, 19.98009, 19.98009, 19.98008, 19.98009, 
    19.98003, 19.98002, 19.97994, 19.97997, 19.97992, 19.97997, 19.97996, 
    19.97992, 19.97996, 19.97986, 19.97993, 19.9798, 19.97987, 19.9798, 
    19.97981, 19.97979, 19.97977, 19.97975, 19.97971, 19.97972, 19.97968, 
    19.98006, 19.98004, 19.98004, 19.98001, 19.98, 19.97996, 19.9799, 
    19.97992, 19.97988, 19.97987, 19.97993, 19.97989, 19.98002, 19.98, 
    19.98001, 19.98006, 19.97992, 19.97999, 19.97985, 19.97989, 19.97978, 
    19.97983, 19.97972, 19.97967, 19.97963, 19.97958, 19.98002, 19.98004, 
    19.98001, 19.97997, 19.97994, 19.97989, 19.97989, 19.97988, 19.97985, 
    19.97983, 19.97987, 19.97983, 19.98, 19.97991, 19.98005, 19.98, 19.97997, 
    19.97999, 19.97992, 19.97991, 19.97985, 19.97988, 19.97968, 19.97977, 
    19.97953, 19.9796, 19.98005, 19.98002, 19.97995, 19.97999, 19.97989, 
    19.97986, 19.97984, 19.97982, 19.97981, 19.9798, 19.97982, 19.9798, 
    19.97989, 19.97985, 19.97996, 19.97993, 19.97994, 19.97996, 19.97992, 
    19.97987, 19.97987, 19.97986, 19.97982, 19.97989, 19.97967, 19.9798, 
    19.98, 19.97996, 19.97996, 19.97997, 19.97986, 19.9799, 19.9798, 
    19.97983, 19.97978, 19.9798, 19.97981, 19.97984, 19.97986, 19.9799, 
    19.97994, 19.97997, 19.97996, 19.97993, 19.97987, 19.97981, 19.97983, 
    19.97979, 19.97989, 19.97985, 19.97987, 19.97982, 19.97992, 19.97984, 
    19.97994, 19.97993, 19.9799, 19.97985, 19.97983, 19.97982, 19.97983, 
    19.97987, 19.97988, 19.9799, 19.97991, 19.97993, 19.97995, 19.97994, 
    19.97992, 19.97987, 19.97982, 19.97977, 19.97976, 19.9797, 19.97975, 
    19.97967, 19.97974, 19.97963, 19.97983, 19.97974, 19.9799, 19.97989, 
    19.97985, 19.97978, 19.97982, 19.97977, 19.97988, 19.97993, 19.97994, 
    19.97997, 19.97994, 19.97994, 19.97992, 19.97993, 19.97987, 19.9799, 
    19.97981, 19.97978, 19.97968, 19.97963, 19.97957, 19.97954, 19.97953, 
    19.97953,
  19.98076, 19.98071, 19.98072, 19.98068, 19.9807, 19.98068, 19.98075, 
    19.98071, 19.98074, 19.98076, 19.9806, 19.98068, 19.98052, 19.98057, 
    19.98044, 19.98052, 19.98042, 19.98044, 19.98038, 19.9804, 19.98033, 
    19.98038, 19.98029, 19.98034, 19.98033, 19.98038, 19.98066, 19.98061, 
    19.98067, 19.98066, 19.98066, 19.9807, 19.98072, 19.98077, 19.98076, 
    19.98073, 19.98066, 19.98068, 19.98062, 19.98062, 19.98055, 19.98058, 
    19.98046, 19.9805, 19.9804, 19.98042, 19.9804, 19.98041, 19.9804, 
    19.98044, 19.98042, 19.98045, 19.98057, 19.98054, 19.98064, 19.98071, 
    19.98075, 19.98078, 19.98078, 19.98077, 19.98073, 19.98069, 19.98066, 
    19.98064, 19.98062, 19.98056, 19.98053, 19.98046, 19.98047, 19.98045, 
    19.98043, 19.98039, 19.9804, 19.98038, 19.98045, 19.9804, 19.98048, 
    19.98046, 19.98061, 19.98067, 19.9807, 19.98072, 19.98078, 19.98074, 
    19.98075, 19.98072, 19.9807, 19.98071, 19.98064, 19.98066, 19.98052, 
    19.98059, 19.98043, 19.98046, 19.98042, 19.98044, 19.9804, 19.98044, 
    19.98038, 19.98036, 19.98037, 19.98034, 19.98044, 19.9804, 19.98071, 
    19.98071, 19.9807, 19.98073, 19.98074, 19.98077, 19.98074, 19.98073, 
    19.98069, 19.98067, 19.98066, 19.98062, 19.98057, 19.98051, 19.98046, 
    19.98043, 19.98045, 19.98043, 19.98045, 19.98046, 19.98037, 19.98042, 
    19.98034, 19.98034, 19.98038, 19.98034, 19.9807, 19.98071, 19.98075, 
    19.98072, 19.98077, 19.98074, 19.98073, 19.98066, 19.98065, 19.98064, 
    19.98061, 19.98058, 19.98052, 19.98047, 19.98042, 19.98043, 19.98043, 
    19.98042, 19.98044, 19.98041, 19.98041, 19.98042, 19.98034, 19.98037, 
    19.98034, 19.98036, 19.98071, 19.98069, 19.9807, 19.98068, 19.9807, 
    19.98064, 19.98063, 19.98055, 19.98058, 19.98053, 19.98057, 19.98057, 
    19.98053, 19.98057, 19.98047, 19.98054, 19.98042, 19.98048, 19.98041, 
    19.98042, 19.9804, 19.98038, 19.98036, 19.98032, 19.98033, 19.98029, 
    19.98067, 19.98064, 19.98065, 19.98062, 19.9806, 19.98057, 19.98051, 
    19.98053, 19.98049, 19.98048, 19.98054, 19.9805, 19.98063, 19.98061, 
    19.98062, 19.98067, 19.98052, 19.9806, 19.98046, 19.9805, 19.98039, 
    19.98044, 19.98033, 19.98029, 19.98024, 19.98019, 19.98063, 19.98065, 
    19.98062, 19.98058, 19.98055, 19.9805, 19.9805, 19.98049, 19.98046, 
    19.98044, 19.98048, 19.98044, 19.9806, 19.98052, 19.98065, 19.98061, 
    19.98058, 19.9806, 19.98053, 19.98052, 19.98046, 19.98049, 19.9803, 
    19.98038, 19.98015, 19.98021, 19.98065, 19.98063, 19.98056, 19.98059, 
    19.9805, 19.98047, 19.98045, 19.98043, 19.98042, 19.98041, 19.98043, 
    19.98041, 19.9805, 19.98046, 19.98057, 19.98054, 19.98055, 19.98057, 
    19.98053, 19.98048, 19.98048, 19.98047, 19.98043, 19.9805, 19.98029, 
    19.98042, 19.98061, 19.98057, 19.98056, 19.98058, 19.98047, 19.98051, 
    19.98041, 19.98044, 19.98039, 19.98042, 19.98042, 19.98045, 19.98046, 
    19.98051, 19.98055, 19.98058, 19.98057, 19.98054, 19.98048, 19.98042, 
    19.98044, 19.9804, 19.9805, 19.98046, 19.98048, 19.98043, 19.98053, 
    19.98045, 19.98055, 19.98054, 19.98051, 19.98046, 19.98044, 19.98043, 
    19.98044, 19.98048, 19.98049, 19.98051, 19.98052, 19.98054, 19.98056, 
    19.98055, 19.98053, 19.98048, 19.98043, 19.98038, 19.98037, 19.98032, 
    19.98036, 19.98029, 19.98035, 19.98024, 19.98044, 19.98035, 19.98051, 
    19.9805, 19.98046, 19.98039, 19.98043, 19.98039, 19.98049, 19.98054, 
    19.98055, 19.98058, 19.98055, 19.98055, 19.98053, 19.98054, 19.98048, 
    19.98051, 19.98042, 19.98039, 19.98029, 19.98024, 19.98018, 19.98016, 
    19.98015, 19.98014,
  19.98279, 19.98275, 19.98276, 19.98272, 19.98274, 19.98271, 19.98278, 
    19.98274, 19.98277, 19.98279, 19.98264, 19.98271, 19.98256, 19.98261, 
    19.98249, 19.98257, 19.98248, 19.98249, 19.98244, 19.98245, 19.98239, 
    19.98243, 19.98235, 19.9824, 19.98239, 19.98243, 19.9827, 19.98265, 
    19.9827, 19.98269, 19.9827, 19.98274, 19.98276, 19.9828, 19.98279, 
    19.98276, 19.98269, 19.98272, 19.98266, 19.98266, 19.98259, 19.98262, 
    19.98251, 19.98254, 19.98245, 19.98248, 19.98245, 19.98246, 19.98245, 
    19.98249, 19.98247, 19.9825, 19.98262, 19.98258, 19.98268, 19.98274, 
    19.98278, 19.98281, 19.98281, 19.9828, 19.98276, 19.98272, 19.98269, 
    19.98268, 19.98266, 19.9826, 19.98257, 19.98251, 19.98252, 19.9825, 
    19.98248, 19.98245, 19.98245, 19.98244, 19.9825, 19.98246, 19.98252, 
    19.98251, 19.98265, 19.98271, 19.98273, 19.98275, 19.9828, 19.98277, 
    19.98278, 19.98275, 19.98273, 19.98274, 19.98268, 19.9827, 19.98257, 
    19.98263, 19.98248, 19.98252, 19.98247, 19.98249, 19.98246, 19.98249, 
    19.98243, 19.98242, 19.98243, 19.9824, 19.98249, 19.98245, 19.98274, 
    19.98274, 19.98273, 19.98277, 19.98277, 19.9828, 19.98277, 19.98276, 
    19.98273, 19.98271, 19.98269, 19.98266, 19.98261, 19.98256, 19.98251, 
    19.98248, 19.9825, 19.98249, 19.9825, 19.98251, 19.98242, 19.98247, 
    19.9824, 19.9824, 19.98244, 19.9824, 19.98274, 19.98275, 19.98278, 
    19.98275, 19.9828, 19.98277, 19.98276, 19.9827, 19.98269, 19.98268, 
    19.98265, 19.98262, 19.98257, 19.98252, 19.98248, 19.98248, 19.98248, 
    19.98247, 19.98249, 19.98247, 19.98246, 19.98247, 19.9824, 19.98242, 
    19.9824, 19.98242, 19.98274, 19.98273, 19.98274, 19.98272, 19.98273, 
    19.98268, 19.98266, 19.98259, 19.98262, 19.98257, 19.98262, 19.98261, 
    19.98257, 19.98261, 19.98252, 19.98258, 19.98247, 19.98253, 19.98247, 
    19.98248, 19.98246, 19.98244, 19.98242, 19.98238, 19.98239, 19.98235, 
    19.9827, 19.98268, 19.98268, 19.98266, 19.98265, 19.98261, 19.98255, 
    19.98257, 19.98254, 19.98253, 19.98259, 19.98255, 19.98267, 19.98265, 
    19.98266, 19.9827, 19.98257, 19.98264, 19.98251, 19.98255, 19.98244, 
    19.9825, 19.98239, 19.98235, 19.98231, 19.98226, 19.98267, 19.98269, 
    19.98266, 19.98262, 19.98259, 19.98255, 19.98254, 19.98253, 19.98251, 
    19.9825, 19.98253, 19.98249, 19.98265, 19.98256, 19.98269, 19.98265, 
    19.98263, 19.98264, 19.98258, 19.98256, 19.98251, 19.98254, 19.98236, 
    19.98244, 19.98222, 19.98228, 19.98269, 19.98267, 19.9826, 19.98264, 
    19.98254, 19.98252, 19.9825, 19.98248, 19.98248, 19.98246, 19.98249, 
    19.98247, 19.98255, 19.98251, 19.98261, 19.98259, 19.9826, 19.98261, 
    19.98257, 19.98253, 19.98253, 19.98252, 19.98248, 19.98254, 19.98235, 
    19.98247, 19.98265, 19.98261, 19.98261, 19.98262, 19.98252, 19.98256, 
    19.98246, 19.98249, 19.98245, 19.98247, 19.98247, 19.9825, 19.98252, 
    19.98256, 19.98259, 19.98262, 19.98261, 19.98258, 19.98253, 19.98248, 
    19.98249, 19.98245, 19.98255, 19.98251, 19.98252, 19.98248, 19.98258, 
    19.9825, 19.9826, 19.98259, 19.98256, 19.98251, 19.98249, 19.98248, 
    19.98249, 19.98253, 19.98253, 19.98256, 19.98257, 19.98259, 19.9826, 
    19.98259, 19.98257, 19.98253, 19.98249, 19.98244, 19.98243, 19.98238, 
    19.98242, 19.98235, 19.98241, 19.9823, 19.98249, 19.98241, 19.98256, 
    19.98254, 19.98251, 19.98245, 19.98248, 19.98244, 19.98253, 19.98258, 
    19.9826, 19.98262, 19.98259, 19.9826, 19.98257, 19.98258, 19.98253, 
    19.98256, 19.98247, 19.98244, 19.98236, 19.9823, 19.98225, 19.98223, 
    19.98222, 19.98222,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7221541, 0.7221522, 0.7221526, 0.7221511, 0.7221519, 0.722151, 0.7221537, 
    0.7221522, 0.7221531, 0.7221539, 0.7221482, 0.722151, 0.7221454, 
    0.7221472, 0.7221427, 0.7221456, 0.7221421, 0.7221428, 0.7221407, 
    0.7221413, 0.7221386, 0.7221404, 0.7221373, 0.7221391, 0.7221388, 
    0.7221405, 0.7221505, 0.7221486, 0.7221506, 0.7221503, 0.7221504, 
    0.7221519, 0.7221527, 0.7221542, 0.7221539, 0.7221528, 0.7221502, 
    0.7221511, 0.7221489, 0.722149, 0.7221465, 0.7221476, 0.7221435, 
    0.7221447, 0.7221413, 0.7221421, 0.7221413, 0.7221416, 0.7221413, 
    0.7221426, 0.722142, 0.7221431, 0.7221474, 0.7221462, 0.7221498, 
    0.7221521, 0.7221536, 0.7221547, 0.7221546, 0.7221543, 0.7221528, 
    0.7221514, 0.7221503, 0.7221497, 0.722149, 0.7221469, 0.7221457, 
    0.7221432, 0.7221437, 0.7221429, 0.7221422, 0.722141, 0.7221412, 
    0.7221407, 0.7221429, 0.7221414, 0.7221439, 0.7221432, 0.7221488, 
    0.7221509, 0.7221518, 0.7221525, 0.7221544, 0.7221531, 0.7221536, 
    0.7221524, 0.7221516, 0.722152, 0.7221496, 0.7221506, 0.7221457, 
    0.7221478, 0.7221423, 0.7221436, 0.722142, 0.7221428, 0.7221414, 
    0.7221426, 0.7221404, 0.72214, 0.7221403, 0.722139, 0.7221428, 0.7221413, 
    0.722152, 0.7221519, 0.7221516, 0.7221529, 0.722153, 0.7221542, 
    0.7221532, 0.7221527, 0.7221516, 0.7221509, 0.7221503, 0.7221488, 
    0.7221473, 0.7221451, 0.7221435, 0.7221425, 0.7221431, 0.7221425, 
    0.7221432, 0.7221435, 0.7221401, 0.722142, 0.7221392, 0.7221394, 
    0.7221406, 0.7221394, 0.7221519, 0.7221523, 0.7221535, 0.7221525, 
    0.7221543, 0.7221534, 0.7221528, 0.7221505, 0.72215, 0.7221496, 
    0.7221487, 0.7221475, 0.7221455, 0.7221438, 0.7221422, 0.7221423, 
    0.7221422, 0.7221419, 0.7221428, 0.7221417, 0.7221416, 0.722142, 
    0.7221394, 0.7221401, 0.7221394, 0.7221398, 0.7221522, 0.7221515, 
    0.7221519, 0.7221513, 0.7221517, 0.7221497, 0.7221492, 0.7221465, 
    0.7221476, 0.7221458, 0.7221474, 0.7221471, 0.7221457, 0.7221473, 
    0.7221438, 0.7221462, 0.7221419, 0.7221442, 0.7221417, 0.7221422, 
    0.7221414, 0.7221407, 0.7221399, 0.7221384, 0.7221388, 0.7221375, 
    0.7221506, 0.7221498, 0.7221499, 0.7221491, 0.7221485, 0.7221472, 
    0.722145, 0.7221458, 0.7221444, 0.7221441, 0.7221463, 0.7221449, 
    0.7221493, 0.7221486, 0.722149, 0.7221506, 0.7221456, 0.7221482, 
    0.7221435, 0.7221448, 0.7221408, 0.7221428, 0.7221389, 0.7221373, 
    0.7221357, 0.7221339, 0.7221494, 0.72215, 0.722149, 0.7221476, 0.7221464, 
    0.7221448, 0.7221446, 0.7221443, 0.7221435, 0.7221428, 0.7221442, 
    0.7221426, 0.7221484, 0.7221454, 0.7221501, 0.7221487, 0.7221477, 
    0.7221482, 0.7221459, 0.7221454, 0.7221432, 0.7221443, 0.7221377, 
    0.7221406, 0.7221324, 0.7221347, 0.7221501, 0.7221494, 0.7221469, 
    0.7221481, 0.7221447, 0.7221438, 0.7221431, 0.7221423, 0.7221422, 
    0.7221416, 0.7221425, 0.7221417, 0.7221448, 0.7221434, 0.7221472, 
    0.7221463, 0.7221467, 0.7221472, 0.7221457, 0.7221442, 0.7221441, 
    0.7221437, 0.7221423, 0.7221447, 0.7221373, 0.7221419, 0.7221486, 
    0.7221472, 0.722147, 0.7221476, 0.7221439, 0.7221453, 0.7221417, 
    0.7221426, 0.722141, 0.7221418, 0.7221419, 0.7221429, 0.7221436, 
    0.7221452, 0.7221465, 0.7221475, 0.7221472, 0.7221462, 0.7221441, 
    0.7221422, 0.7221426, 0.7221411, 0.7221449, 0.7221434, 0.7221439, 
    0.7221423, 0.7221459, 0.7221429, 0.7221466, 0.7221463, 0.7221453, 
    0.7221432, 0.7221428, 0.7221423, 0.7221426, 0.722144, 0.7221442, 
    0.7221453, 0.7221456, 0.7221463, 0.722147, 0.7221464, 0.7221458, 
    0.722144, 0.7221425, 0.7221407, 0.7221403, 0.7221383, 0.72214, 0.7221373, 
    0.7221395, 0.7221356, 0.7221427, 0.7221396, 0.7221452, 0.7221446, 
    0.7221435, 0.722141, 0.7221424, 0.7221408, 0.7221443, 0.7221461, 
    0.7221466, 0.7221474, 0.7221465, 0.7221466, 0.7221457, 0.722146, 
    0.7221439, 0.7221451, 0.7221419, 0.7221408, 0.7221376, 0.7221356, 
    0.7221336, 0.7221327, 0.7221324, 0.7221323 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  1.027984e-20, -3.597945e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -2.055969e-20, 1.027984e-20, -2.055969e-20, 
    1.027984e-20, 1.541976e-20, -2.006177e-36, 0, 5.139921e-21, 
    -4.111937e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    2.006177e-36, -2.006177e-36, -1.541976e-20, -5.139921e-21, 5.139921e-20, 
    -2.569961e-20, 0, 1.541976e-20, 1.027984e-20, 1.541976e-20, 1.027984e-20, 
    5.139921e-21, 5.139921e-20, -1.027984e-20, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, -4.111937e-20, -2.569961e-20, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-20, 2.055969e-20, 1.027984e-20, 
    1.027984e-20, -3.597945e-20, 0, 0, 1.027984e-20, -5.653913e-20, 
    -1.027984e-20, -1.541976e-20, 2.569961e-20, -1.541976e-20, 5.139921e-21, 
    -1.027984e-20, -4.111937e-20, 5.139921e-21, 1.541976e-20, -2.569961e-20, 
    1.541976e-20, -2.055969e-20, -2.006177e-36, 2.569961e-20, -2.569961e-20, 
    -3.083953e-20, -2.055969e-20, -3.597945e-20, -4.111937e-20, 3.083953e-20, 
    1.541976e-20, -3.597945e-20, 1.541976e-20, 2.055969e-20, 1.027984e-20, 
    -2.569961e-20, -1.027984e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, 2.569961e-20, 5.139921e-21, -5.139921e-21, 2.569961e-20, 
    -2.055969e-20, -1.541976e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    4.625929e-20, 2.569961e-20, -2.569961e-20, -2.569961e-20, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, -2.055969e-20, -1.541976e-20, 
    2.569961e-20, -2.569961e-20, -5.139921e-21, -2.055969e-20, 2.055969e-20, 
    2.006177e-36, 3.083953e-20, -2.055969e-20, -1.541976e-20, -4.111937e-20, 
    2.006177e-36, 1.541976e-20, 0, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, 2.006177e-36, 
    3.597945e-20, -3.083953e-20, 5.139921e-21, -3.597945e-20, -1.027984e-20, 
    -1.027984e-20, 2.569961e-20, 0, 0, -2.055969e-20, 1.541976e-20, 
    1.027984e-20, 1.027984e-20, 2.569961e-20, 3.083953e-20, 5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, 2.569961e-20, 2.055969e-20, 
    -5.139921e-21, 2.569961e-20, 2.569961e-20, 3.597945e-20, -3.083953e-20, 
    0, -5.139921e-21, 5.139921e-21, 0, -1.027984e-20, 3.597945e-20, 
    -5.139921e-21, -2.006177e-36, -5.139921e-21, -1.541976e-20, 2.055969e-20, 
    -2.569961e-20, -1.541976e-20, 2.055969e-20, 1.541976e-20, -1.541976e-20, 
    2.569961e-20, -5.139921e-21, -2.055969e-20, 2.055969e-20, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, -1.027984e-20, -2.006177e-36, -4.111937e-20, 
    1.541976e-20, -5.139921e-21, 2.569961e-20, -1.027984e-20, 2.055969e-20, 
    -2.569961e-20, 2.569961e-20, 5.139921e-21, -1.027984e-20, 0, 
    4.625929e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 2.055969e-20, 
    1.027984e-20, 1.541976e-20, 1.541976e-20, 4.625929e-20, 5.139921e-21, 
    -2.055969e-20, 3.597945e-20, 5.139921e-21, 2.569961e-20, 2.569961e-20, 0, 
    -2.569961e-20, 1.027984e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    2.055969e-20, 2.055969e-20, 2.569961e-20, 2.569961e-20, -1.027984e-20, 
    -2.006177e-36, -2.055969e-20, 2.055969e-20, -1.541976e-20, -2.055969e-20, 
    2.055969e-20, 2.569961e-20, 1.027984e-20, -1.027984e-20, 2.006177e-36, 
    -2.055969e-20, -1.027984e-20, 5.139921e-21, 2.055969e-20, 1.027984e-20, 
    -3.083953e-20, 0, 0, -3.597945e-20, 1.541976e-20, 3.083953e-20, 
    2.569961e-20, -3.597945e-20, -2.006177e-36, 1.541976e-20, -1.027984e-20, 
    3.083953e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    2.569961e-20, 1.027984e-20, -2.569961e-20, 2.569961e-20, -1.027984e-20, 
    1.541976e-20, -2.055969e-20, 5.139921e-21, 1.027984e-20, -3.083953e-20, 
    -5.139921e-21, 5.139921e-21, 2.055969e-20, -3.597945e-20, -5.139921e-21, 
    5.139921e-21, 2.055969e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    2.569961e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, -1.027984e-20, 
    1.027984e-20, -1.541976e-20, 2.569961e-20, 1.541976e-20, 5.139921e-21, 
    -1.027984e-20, 1.541976e-20, -2.569961e-20, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -2.055969e-20, 1.541976e-20, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, -2.006177e-36, -1.027984e-20, -1.027984e-20, 
    -1.541976e-20, 2.055969e-20, -2.006177e-36, -5.139921e-21, -2.569961e-20, 
    2.006177e-36, 5.139921e-21, 1.027984e-20, 1.027984e-20, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, 2.006177e-36, -2.569961e-20, -1.027984e-20, 
    -1.027984e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, -3.083953e-20, 
    1.541976e-20, 1.541976e-20, 1.541976e-20, 5.139921e-21, 1.541976e-20, 
    -2.569961e-20, -2.569961e-20, 1.541976e-20, -5.139921e-21, -2.569961e-20, 
    0, -5.139921e-21, -5.139921e-21, 1.541976e-20, 2.055969e-20, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 2.569961e-20, 
    2.006177e-36, -1.027984e-20, -2.055969e-20, -2.055969e-20, 5.139921e-21, 
    -2.006177e-36, 1.027984e-20,
  5.139921e-21, -2.569961e-20, 1.541976e-20, 2.055969e-20, 1.541976e-20, 
    -5.139921e-21, -2.569961e-20, -2.055969e-20, -2.569961e-20, 0, 
    -2.569961e-20, -1.541976e-20, 1.541976e-20, 1.541976e-20, 1.541976e-20, 
    3.083953e-20, -5.139921e-21, 0, 2.006177e-36, 2.569961e-20, 0, 
    -5.139921e-21, 0, 5.139921e-21, 5.139921e-21, -1.541976e-20, 
    2.055969e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 
    -2.569961e-20, 0, -2.006177e-36, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, 2.055969e-20, 5.139921e-21, -1.027984e-20, 3.083953e-20, 
    5.139921e-21, 2.569961e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, 
    5.139921e-21, -1.541976e-20, 3.083953e-20, -1.541976e-20, 1.541976e-20, 
    5.139921e-21, -3.597945e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 2.055969e-20, 
    1.027984e-20, -3.597945e-20, 5.139921e-21, 2.055969e-20, 2.055969e-20, 
    -5.139921e-21, 0, 5.139921e-21, -1.541976e-20, 3.597945e-20, 
    -1.541976e-20, 2.055969e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -2.055969e-20, -5.139921e-21, -2.055969e-20, 
    -1.541976e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 0, -1.027984e-20, 2.006177e-36, 
    -2.569961e-20, -5.139921e-21, -5.139921e-21, -2.569961e-20, 
    -2.055969e-20, 2.006177e-36, 5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -2.569961e-20, 2.569961e-20, 1.541976e-20, -1.541976e-20, 0, 
    5.139921e-21, 3.083953e-20, -2.569961e-20, -5.139921e-21, -5.139921e-21, 
    2.055969e-20, 5.139921e-21, 3.083953e-20, 2.569961e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -2.569961e-20, -1.027984e-20, 1.541976e-20, 
    2.569961e-20, -1.541976e-20, -5.139921e-21, -1.027984e-20, -2.055969e-20, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, -1.541976e-20, 0, 
    -2.569961e-20, 1.541976e-20, 1.027984e-20, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -2.055969e-20, -1.541976e-20, 1.027984e-20, 
    2.006177e-36, 0, 1.541976e-20, -5.139921e-21, -1.027984e-20, 0, 
    1.541976e-20, -1.541976e-20, -1.027984e-20, 0, 2.055969e-20, 
    -1.027984e-20, -1.541976e-20, -1.027984e-20, 1.541976e-20, 3.083953e-20, 
    0, 0, 5.139921e-21, 5.139921e-21, -1.541976e-20, -2.055969e-20, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, -2.569961e-20, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, -2.569961e-20, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, 2.055969e-20, 3.083953e-20, 0, 
    -1.027984e-20, 0, 1.027984e-20, -5.139921e-21, -2.569961e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    3.083953e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 2.055969e-20, 
    -5.139921e-21, -1.541976e-20, -1.541976e-20, 1.541976e-20, 2.055969e-20, 
    -1.541976e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, 3.597945e-20, 
    -1.541976e-20, -5.139921e-21, -2.569961e-20, -1.541976e-20, 
    -1.027984e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, 1.027984e-20, 0, -1.027984e-20, 1.541976e-20, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 2.055969e-20, 
    1.027984e-20, -2.055969e-20, -1.541976e-20, 1.027984e-20, 2.569961e-20, 
    -2.055969e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, -2.006177e-36, 
    0, -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    2.569961e-20, 1.027984e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 
    2.569961e-20, -1.027984e-20, -2.055969e-20, 2.569961e-20, 1.027984e-20, 
    2.055969e-20, -1.541976e-20, 3.083953e-20, -2.055969e-20, -1.027984e-20, 
    2.006177e-36, -1.027984e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, -1.541976e-20, 0, 
    -1.027984e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, -1.027984e-20, 2.569961e-20, 
    -2.569961e-20, -1.027984e-20, 1.027984e-20, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, -2.055969e-20, -1.027984e-20, 
    -5.139921e-21, 2.055969e-20, -2.055969e-20, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 1.541976e-20, -2.569961e-20, -2.055969e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -2.055969e-20, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 0, -1.027984e-20, -5.139921e-21, 
    -2.055969e-20, 1.541976e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    3.083953e-20, 1.541976e-20, 5.139921e-21, 3.597945e-20, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, -1.027984e-20, -2.055969e-20, -5.139921e-21, 
    0, 0, -1.027984e-20, 2.055969e-20, 5.139921e-21, -2.055969e-20, 
    -1.027984e-20, 2.006177e-36, 5.139921e-21, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -2.569961e-20, -1.541976e-20,
  3.597945e-20, -2.569961e-20, 1.027984e-20, -2.055969e-20, -1.541976e-20, 
    1.027984e-20, 0, 2.569961e-20, -1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, 3.083953e-20, -5.139921e-21, 
    3.083953e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, 1.027984e-20, 
    -1.027984e-20, -1.027984e-20, 0, -3.083953e-20, -2.569961e-20, 
    5.139921e-21, 2.055969e-20, 1.027984e-20, -2.006177e-36, 2.006177e-36, 
    5.139921e-21, 2.006177e-36, -5.139921e-21, 1.541976e-20, 1.541976e-20, 
    5.139921e-21, -3.083953e-20, 0, 5.139921e-21, -5.139921e-21, 
    1.541976e-20, 5.139921e-21, 2.569961e-20, -1.541976e-20, 2.055969e-20, 
    1.027984e-20, 4.111937e-20, 1.027984e-20, 2.055969e-20, 2.055969e-20, 
    1.541976e-20, -1.541976e-20, 2.569961e-20, 2.006177e-36, 1.027984e-20, 
    5.139921e-21, 1.541976e-20, -2.055969e-20, -2.055969e-20, -2.006177e-36, 
    1.541976e-20, 5.139921e-21, 2.006177e-36, -2.006177e-36, -2.055969e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -2.055969e-20, -2.569961e-20, -1.541976e-20, 3.597945e-20, -1.027984e-20, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, 2.569961e-20, -5.139921e-21, 
    -5.139921e-21, 2.569961e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -2.569961e-20, 1.541976e-20, -2.569961e-20, 5.139921e-21, 5.139921e-21, 
    -4.111937e-20, 5.139921e-21, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    1.027984e-20, -5.139921e-21, -1.541976e-20, -3.597945e-20, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 3.083953e-20, -1.541976e-20, 5.139921e-21, 
    1.027984e-20, 2.055969e-20, -3.083953e-20, -1.541976e-20, -2.569961e-20, 
    -2.055969e-20, 1.541976e-20, 0, 1.541976e-20, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, 1.541976e-20, 2.055969e-20, 
    2.569961e-20, 3.083953e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, -4.111937e-20, 1.027984e-20, -1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, -5.139921e-21, 
    -2.055969e-20, 2.055969e-20, -3.597945e-20, 1.027984e-20, 0, 
    5.139921e-21, -2.569961e-20, -3.597945e-20, 1.541976e-20, -1.541976e-20, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, -2.055969e-20, 
    -5.139921e-21, 3.083953e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, 
    -3.083953e-20, -2.055969e-20, -2.055969e-20, -2.006177e-36, 
    -5.139921e-21, 0, -1.027984e-20, -5.139921e-21, 2.055969e-20, 
    5.139921e-21, -3.083953e-20, 0, -2.569961e-20, 5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 1.027984e-20, 0, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 0, -1.541976e-20, -1.027984e-20, 
    -2.055969e-20, 0, 1.027984e-20, 0, -1.541976e-20, -1.027984e-20, 
    -2.055969e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 1.027984e-20, 
    2.006177e-36, -1.541976e-20, -2.569961e-20, 1.541976e-20, 1.027984e-20, 
    -1.541976e-20, -2.055969e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    1.541976e-20, -5.139921e-21, 5.139921e-21, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 2.006177e-36, -2.055969e-20, 5.139921e-21, 0, 
    -2.006177e-36, 1.541976e-20, -1.027984e-20, 0, 1.541976e-20, 
    -5.139921e-21, 2.055969e-20, 2.055969e-20, 0, 2.055969e-20, 
    -2.055969e-20, -1.541976e-20, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -2.006177e-36, 5.139921e-21, 1.027984e-20, -2.569961e-20, -1.027984e-20, 
    2.055969e-20, 5.139921e-21, -5.139921e-21, -2.055969e-20, 2.055969e-20, 
    1.027984e-20, 2.055969e-20, 1.541976e-20, 1.027984e-20, -2.006177e-36, 
    -1.541976e-20, -1.541976e-20, 1.541976e-20, 1.027984e-20, 3.597945e-20, 
    1.541976e-20, 2.055969e-20, 3.083953e-20, 2.055969e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-20, 1.541976e-20, -1.541976e-20, 
    5.139921e-21, 3.083953e-20, -1.541976e-20, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, 2.006177e-36, -2.055969e-20, -2.055969e-20, -3.083953e-20, 
    -3.597945e-20, -5.139921e-21, -1.541976e-20, 3.597945e-20, 1.027984e-20, 
    3.083953e-20, -2.055969e-20, -1.541976e-20, 3.083953e-20, 1.541976e-20, 
    -1.027984e-20, 2.569961e-20, -2.055969e-20, -1.541976e-20, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 0, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, 1.541976e-20, 
    2.055969e-20, -1.541976e-20, -1.027984e-20, 1.027984e-20, 2.055969e-20, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, 1.027984e-20, 
    1.541976e-20, 2.569961e-20, -1.027984e-20, -1.027984e-20, 2.055969e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-20, 1.027984e-20, 1.541976e-20, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, 3.083953e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -2.055969e-20, 5.139921e-21, 0, 
    -1.541976e-20, -5.139921e-21, -2.055969e-20, 5.139921e-21, 2.055969e-20, 
    3.083953e-20, 3.597945e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    2.055969e-20, 1.027984e-20, 0, 2.569961e-20,
  -2.055969e-20, 0, -1.027984e-20, 1.541976e-20, -1.027984e-20, 5.139921e-21, 
    2.569961e-20, 1.027984e-20, 1.541976e-20, -3.597945e-20, 0, 2.055969e-20, 
    -5.139921e-21, 5.139921e-21, 2.055969e-20, 4.625929e-20, 2.055969e-20, 
    3.597945e-20, 2.006177e-36, -5.139921e-21, 1.027984e-20, 1.541976e-20, 
    2.055969e-20, 0, 2.055969e-20, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, 1.027984e-20, -3.597945e-20, 3.597945e-20, 2.055969e-20, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, -1.027984e-20, -4.625929e-20, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -5.139921e-20, -1.027984e-20, -3.597945e-20, -5.139921e-21, 5.139921e-21, 
    4.625929e-20, -5.139921e-21, 2.055969e-20, -2.055969e-20, -2.055969e-20, 
    -2.569961e-20, 1.027984e-20, 2.055969e-20, 1.027984e-20, 2.055969e-20, 0, 
    3.083953e-20, 3.083953e-20, 1.541976e-20, 2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 2.569961e-20, -2.569961e-20, -2.569961e-20, 1.027984e-20, 
    2.006177e-36, -4.111937e-20, -1.027984e-20, -1.541976e-20, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, 3.083953e-20, -2.055969e-20, -1.541976e-20, 
    2.055969e-20, 5.139921e-21, 2.006177e-36, -5.139921e-21, -3.597945e-20, 
    3.083953e-20, 5.139921e-21, 4.111937e-20, -2.006177e-36, 1.541976e-20, 
    3.083953e-20, 1.027984e-20, 0, 2.006177e-36, 5.139921e-21, -5.139921e-21, 
    -2.055969e-20, 1.541976e-20, -5.139921e-21, 5.139921e-21, -1.541976e-20, 
    1.541976e-20, -5.139921e-21, 2.569961e-20, 1.541976e-20, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, -1.541976e-20, -3.597945e-20, -2.055969e-20, 
    1.027984e-20, -2.569961e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    2.006177e-36, -2.055969e-20, -2.569961e-20, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, -2.055969e-20, 
    5.139921e-21, -1.027984e-20, -2.006177e-36, 0, 5.139921e-21, 
    1.541976e-20, 1.541976e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 3.083953e-20, -2.006177e-36, -5.139921e-21, -2.569961e-20, 
    5.139921e-21, 2.569961e-20, 0, -1.027984e-20, 1.027984e-20, 
    -1.027984e-20, -2.055969e-20, 1.027984e-20, 0, -1.541976e-20, 
    -2.006177e-36, 0, 1.541976e-20, -1.027984e-20, -2.006177e-36, 
    2.569961e-20, -3.083953e-20, 1.541976e-20, -5.139921e-21, -2.055969e-20, 
    -2.569961e-20, 1.027984e-20, -5.139921e-21, -1.541976e-20, 1.541976e-20, 
    3.597945e-20, -2.055969e-20, 2.055969e-20, 0, -5.139921e-21, 
    -1.541976e-20, 2.055969e-20, 5.139921e-21, 0, 1.027984e-20, 
    -5.139921e-21, -3.597945e-20, 5.139921e-21, 1.027984e-20, 0, 
    1.027984e-20, -3.597945e-20, 1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -2.055969e-20, -1.027984e-20, 0, 
    2.055969e-20, 1.541976e-20, 0, 3.083953e-20, -1.027984e-20, 
    -1.027984e-20, -2.055969e-20, 0, -2.569961e-20, -5.139921e-21, 
    5.139921e-21, 2.569961e-20, -1.027984e-20, 4.111937e-20, -1.027984e-20, 
    1.027984e-20, -6.167906e-20, 5.139921e-21, 1.541976e-20, 2.055969e-20, 
    -2.055969e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 2.569961e-20, 
    0, 2.055969e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 2.006177e-36, 
    -2.055969e-20, 5.139921e-21, -3.597945e-20, 1.541976e-20, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -2.569961e-20, -3.083953e-20, 
    1.541976e-20, -2.055969e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, -1.541976e-20, 2.569961e-20, -2.569961e-20, -5.139921e-21, 
    1.541976e-20, 2.569961e-20, 1.027984e-20, 1.027984e-20, 2.569961e-20, 
    2.055969e-20, 2.055969e-20, 4.111937e-20, 2.055969e-20, -1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 5.139921e-21, 3.083953e-20, 1.541976e-20, 
    1.541976e-20, -1.541976e-20, 2.569961e-20, 1.027984e-20, 0, 4.111937e-20, 
    5.139921e-21, 1.541976e-20, -2.055969e-20, -2.569961e-20, 4.111937e-20, 
    2.006177e-36, 5.139921e-21, 1.027984e-20, -1.027984e-20, 0, 
    -1.027984e-20, 5.139921e-21, -1.027984e-20, -1.027984e-20, -1.027984e-20, 
    1.541976e-20, 1.541976e-20, -4.625929e-20, 2.569961e-20, -3.597945e-20, 
    -2.569961e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, -3.597945e-20, 
    -3.083953e-20, 1.541976e-20, -2.055969e-20, -3.597945e-20, -2.055969e-20, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, -5.139921e-21, 3.597945e-20, 
    0, 2.006177e-36, -2.569961e-20, 5.139921e-21, 2.055969e-20, 
    -2.569961e-20, 1.541976e-20, -3.083953e-20, -2.055969e-20, 0, 
    -2.055969e-20, 0, 3.083953e-20, -2.006177e-36, 3.083953e-20, 
    3.083953e-20, 3.083953e-20, -3.597945e-20, 5.139921e-21, 0, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, -1.541976e-20, -2.055969e-20, 
    5.139921e-21, 4.625929e-20, 2.006177e-36, -2.006177e-36, 0, 
    -1.541976e-20, -2.055969e-20,
  -2.569961e-20, -1.027984e-20, 2.569961e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -1.027984e-20, -1.541976e-20, -1.541976e-20, 5.139921e-21, 0, 
    5.139921e-21, -1.027984e-20, 2.569961e-20, -2.055969e-20, -2.055969e-20, 
    1.541976e-20, 2.055969e-20, 5.139921e-21, -1.541976e-20, 1.027984e-20, 
    -1.027984e-20, 2.055969e-20, -3.597945e-20, 2.055969e-20, 5.139921e-21, 
    -2.569961e-20, -5.139921e-21, 4.625929e-20, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 3.597945e-20, 
    -3.597945e-20, 1.541976e-20, -2.569961e-20, 5.139921e-21, -2.055969e-20, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, 0, 0, -1.027984e-20, 
    2.569961e-20, 2.006177e-36, 5.139921e-21, -3.083953e-20, -2.569961e-20, 
    2.569961e-20, 5.139921e-21, -2.569961e-20, 1.027984e-20, 2.055969e-20, 
    2.055969e-20, -3.083953e-20, 4.111937e-20, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -2.569961e-20, -1.541976e-20, -3.597945e-20, 1.541976e-20, 
    -1.541976e-20, 2.006177e-36, -2.569961e-20, 1.027984e-20, -3.083953e-20, 
    -2.055969e-20, 1.027984e-20, -1.541976e-20, 0, 5.139921e-21, 
    5.139921e-21, -3.083953e-20, -2.569961e-20, 3.597945e-20, -2.569961e-20, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, 2.006177e-36, -2.006177e-36, 
    -1.027984e-20, -3.597945e-20, 5.139921e-21, -1.541976e-20, 2.055969e-20, 
    2.055969e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, -2.055969e-20, 
    -3.083953e-20, 2.055969e-20, -1.541976e-20, 1.027984e-20, 2.055969e-20, 
    2.006177e-36, 0, 0, 3.083953e-20, 0, 1.541976e-20, -2.569961e-20, 
    2.055969e-20, -1.027984e-20, -1.541976e-20, -2.055969e-20, -3.083953e-20, 
    -1.027984e-20, 4.111937e-20, 1.541976e-20, -2.006177e-36, 2.055969e-20, 
    -2.055969e-20, -1.541976e-20, -5.139921e-21, 2.055969e-20, -1.541976e-20, 
    -1.541976e-20, -1.541976e-20, 1.027984e-20, 1.027984e-20, -2.055969e-20, 
    0, 2.569961e-20, -5.139921e-21, 2.055969e-20, 2.055969e-20, 
    -4.111937e-20, 2.569961e-20, 1.027984e-20, -1.541976e-20, 2.006177e-36, 
    -1.541976e-20, -2.006177e-36, -2.055969e-20, -2.055969e-20, 5.139921e-21, 
    -2.055969e-20, 3.597945e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, -1.541976e-20, 
    5.139921e-21, -2.055969e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, 2.055969e-20, -2.569961e-20, 2.055969e-20, -3.597945e-20, 
    -2.569961e-20, 5.139921e-21, 1.541976e-20, 3.083953e-20, -1.541976e-20, 
    2.055969e-20, 4.111937e-20, 2.055969e-20, 0, 1.541976e-20, 1.027984e-20, 
    5.139921e-21, 1.027984e-20, 1.541976e-20, 5.139921e-21, 2.006177e-36, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 2.055969e-20, 2.569961e-20, 5.139921e-21, 
    -1.541976e-20, 1.541976e-20, 1.541976e-20, -2.569961e-20, 2.006177e-36, 
    2.569961e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 2.006177e-36, -1.541976e-20, 
    3.083953e-20, 5.139921e-21, 2.055969e-20, 3.083953e-20, 1.541976e-20, 
    -4.111937e-20, -1.027984e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, 
    0, 2.055969e-20, 2.006177e-36, 5.139921e-21, 1.541976e-20, -2.569961e-20, 
    1.027984e-20, -3.083953e-20, 1.541976e-20, 2.569961e-20, -5.139921e-21, 
    -5.139921e-21, 3.083953e-20, -5.139921e-21, 5.139921e-21, -3.597945e-20, 
    -1.541976e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, -2.055969e-20, 
    1.027984e-20, -2.006177e-36, 1.541976e-20, -2.055969e-20, -1.541976e-20, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, -2.006177e-36, 
    -5.139921e-21, 0, -5.139921e-21, -2.055969e-20, -5.139921e-21, 
    -2.055969e-20, -2.055969e-20, 1.027984e-20, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, 2.055969e-20, -1.541976e-20, -3.083953e-20, -5.139921e-21, 
    1.027984e-20, -5.139921e-21, 3.083953e-20, 0, 2.055969e-20, 
    -3.083953e-20, 2.006177e-36, -1.541976e-20, -2.569961e-20, -1.027984e-20, 
    5.139921e-21, 2.055969e-20, -2.569961e-20, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 2.055969e-20, -5.139921e-21, -1.541976e-20, 
    -2.055969e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, -2.055969e-20, 
    1.027984e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 2.006177e-36, 
    5.139921e-21, 0, -1.027984e-20, -2.006177e-36, -4.111937e-20, 
    1.541976e-20, 2.055969e-20, 2.569961e-20, 2.569961e-20, -1.027984e-20, 0, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, -3.083953e-20, 2.055969e-20, 
    -1.541976e-20, 2.055969e-20, -2.055969e-20, -1.541976e-20, 2.569961e-20, 
    -3.597945e-20, -1.541976e-20, 1.541976e-20, -1.027984e-20, 1.541976e-20, 
    -2.055969e-20, 0, -2.055969e-20, -2.006177e-36, 0, 5.139921e-21, 
    2.006177e-36, -1.027984e-20, -1.541976e-20, 1.541976e-20, -2.006177e-36, 
    2.006177e-36, 1.027984e-20,
  8.597411e-29, 8.59739e-29, 8.597394e-29, 8.597377e-29, 8.597387e-29, 
    8.597376e-29, 8.597407e-29, 8.597389e-29, 8.597401e-29, 8.597409e-29, 
    8.597345e-29, 8.597377e-29, 8.597312e-29, 8.597332e-29, 8.597281e-29, 
    8.597315e-29, 8.597274e-29, 8.597282e-29, 8.597258e-29, 8.597265e-29, 
    8.597235e-29, 8.597255e-29, 8.597219e-29, 8.59724e-29, 8.597236e-29, 
    8.597256e-29, 8.59737e-29, 8.597349e-29, 8.597372e-29, 8.597368e-29, 
    8.59737e-29, 8.597386e-29, 8.597395e-29, 8.597413e-29, 8.597409e-29, 
    8.597396e-29, 8.597367e-29, 8.597377e-29, 8.597352e-29, 8.597352e-29, 
    8.597324e-29, 8.597337e-29, 8.59729e-29, 8.597303e-29, 8.597265e-29, 
    8.597274e-29, 8.597265e-29, 8.597268e-29, 8.597265e-29, 8.59728e-29, 
    8.597273e-29, 8.597286e-29, 8.597334e-29, 8.597321e-29, 8.597363e-29, 
    8.597389e-29, 8.597406e-29, 8.597418e-29, 8.597416e-29, 8.597413e-29, 
    8.597396e-29, 8.597381e-29, 8.597369e-29, 8.59736e-29, 8.597352e-29, 
    8.597328e-29, 8.597316e-29, 8.597287e-29, 8.597292e-29, 8.597284e-29, 
    8.597275e-29, 8.597262e-29, 8.597264e-29, 8.597257e-29, 8.597284e-29, 
    8.597266e-29, 8.597295e-29, 8.597287e-29, 8.59735e-29, 8.597374e-29, 
    8.597384e-29, 8.597393e-29, 8.597415e-29, 8.5974e-29, 8.597406e-29, 
    8.597392e-29, 8.597383e-29, 8.597387e-29, 8.59736e-29, 8.597371e-29, 
    8.597315e-29, 8.597339e-29, 8.597277e-29, 8.597292e-29, 8.597273e-29, 
    8.597282e-29, 8.597266e-29, 8.597281e-29, 8.597256e-29, 8.59725e-29, 
    8.597254e-29, 8.597239e-29, 8.597281e-29, 8.597265e-29, 8.597387e-29, 
    8.597387e-29, 8.597384e-29, 8.597398e-29, 8.597399e-29, 8.597413e-29, 
    8.597401e-29, 8.597395e-29, 8.597383e-29, 8.597375e-29, 8.597368e-29, 
    8.597351e-29, 8.597334e-29, 8.597309e-29, 8.59729e-29, 8.597278e-29, 
    8.597286e-29, 8.597279e-29, 8.597286e-29, 8.59729e-29, 8.597252e-29, 
    8.597273e-29, 8.597241e-29, 8.597243e-29, 8.597257e-29, 8.597243e-29, 
    8.597386e-29, 8.59739e-29, 8.597405e-29, 8.597393e-29, 8.597414e-29, 
    8.597402e-29, 8.597396e-29, 8.597371e-29, 8.597365e-29, 8.59736e-29, 
    8.597349e-29, 8.597336e-29, 8.597313e-29, 8.597293e-29, 8.597275e-29, 
    8.597276e-29, 8.597276e-29, 8.597272e-29, 8.597282e-29, 8.59727e-29, 
    8.597268e-29, 8.597273e-29, 8.597243e-29, 8.597252e-29, 8.597243e-29, 
    8.597248e-29, 8.597389e-29, 8.597382e-29, 8.597386e-29, 8.597379e-29, 
    8.597384e-29, 8.597362e-29, 8.597355e-29, 8.597324e-29, 8.597337e-29, 
    8.597316e-29, 8.597334e-29, 8.597331e-29, 8.597316e-29, 8.597334e-29, 
    8.597294e-29, 8.597321e-29, 8.597272e-29, 8.597298e-29, 8.59727e-29, 
    8.597275e-29, 8.597266e-29, 8.597259e-29, 8.59725e-29, 8.597232e-29, 
    8.597236e-29, 8.597221e-29, 8.597372e-29, 8.597363e-29, 8.597363e-29, 
    8.597354e-29, 8.597347e-29, 8.597332e-29, 8.597307e-29, 8.597317e-29, 
    8.5973e-29, 8.597297e-29, 8.597322e-29, 8.597307e-29, 8.597357e-29, 
    8.597349e-29, 8.597354e-29, 8.597371e-29, 8.597315e-29, 8.597343e-29, 
    8.59729e-29, 8.597306e-29, 8.59726e-29, 8.597283e-29, 8.597238e-29, 
    8.597219e-29, 8.597201e-29, 8.59718e-29, 8.597358e-29, 8.597364e-29, 
    8.597353e-29, 8.597338e-29, 8.597324e-29, 8.597305e-29, 8.597303e-29, 
    8.5973e-29, 8.59729e-29, 8.597283e-29, 8.597298e-29, 8.597281e-29, 
    8.597346e-29, 8.597312e-29, 8.597366e-29, 8.59735e-29, 8.597339e-29, 
    8.597343e-29, 8.597318e-29, 8.597312e-29, 8.597287e-29, 8.5973e-29, 
    8.597224e-29, 8.597257e-29, 8.597163e-29, 8.59719e-29, 8.597366e-29, 
    8.597358e-29, 8.597329e-29, 8.597343e-29, 8.597304e-29, 8.597294e-29, 
    8.597286e-29, 8.597276e-29, 8.597275e-29, 8.597269e-29, 8.597279e-29, 
    8.597269e-29, 8.597305e-29, 8.597289e-29, 8.597333e-29, 8.597322e-29, 
    8.597327e-29, 8.597332e-29, 8.597316e-29, 8.597298e-29, 8.597298e-29, 
    8.597292e-29, 8.597276e-29, 8.597304e-29, 8.597219e-29, 8.597271e-29, 
    8.597349e-29, 8.597333e-29, 8.597331e-29, 8.597337e-29, 8.597295e-29, 
    8.59731e-29, 8.597269e-29, 8.59728e-29, 8.597262e-29, 8.597271e-29, 
    8.597272e-29, 8.597284e-29, 8.597291e-29, 8.597309e-29, 8.597324e-29, 
    8.597336e-29, 8.597333e-29, 8.597321e-29, 8.597297e-29, 8.597275e-29, 
    8.59728e-29, 8.597263e-29, 8.597307e-29, 8.597289e-29, 8.597295e-29, 
    8.597277e-29, 8.597317e-29, 8.597283e-29, 8.597325e-29, 8.597322e-29, 
    8.59731e-29, 8.597287e-29, 8.597282e-29, 8.597277e-29, 8.59728e-29, 
    8.597297e-29, 8.597299e-29, 8.597311e-29, 8.597314e-29, 8.597323e-29, 
    8.59733e-29, 8.597324e-29, 8.597316e-29, 8.597297e-29, 8.597278e-29, 
    8.597259e-29, 8.597254e-29, 8.597231e-29, 8.59725e-29, 8.597219e-29, 
    8.597245e-29, 8.5972e-29, 8.597281e-29, 8.597246e-29, 8.59731e-29, 
    8.597303e-29, 8.59729e-29, 8.597262e-29, 8.597277e-29, 8.597259e-29, 
    8.597299e-29, 8.59732e-29, 8.597325e-29, 8.597335e-29, 8.597325e-29, 
    8.597326e-29, 8.597316e-29, 8.597319e-29, 8.597296e-29, 8.597309e-29, 
    8.597272e-29, 8.597259e-29, 8.597222e-29, 8.5972e-29, 8.597177e-29, 
    8.597167e-29, 8.597163e-29, 8.597162e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.397015e-08, 1.400838e-08, 1.400095e-08, 1.403177e-08, 1.401468e-08, 
    1.403486e-08, 1.39779e-08, 1.400989e-08, 1.398947e-08, 1.397359e-08, 
    1.409157e-08, 1.403315e-08, 1.415225e-08, 1.411501e-08, 1.420855e-08, 
    1.414645e-08, 1.422107e-08, 1.420676e-08, 1.424983e-08, 1.423749e-08, 
    1.429254e-08, 1.425552e-08, 1.432108e-08, 1.428371e-08, 1.428955e-08, 
    1.42543e-08, 1.404491e-08, 1.408429e-08, 1.404258e-08, 1.404819e-08, 
    1.404567e-08, 1.401503e-08, 1.399958e-08, 1.396723e-08, 1.397311e-08, 
    1.399686e-08, 1.405072e-08, 1.403245e-08, 1.407851e-08, 1.407747e-08, 
    1.412873e-08, 1.410562e-08, 1.419176e-08, 1.416729e-08, 1.423801e-08, 
    1.422022e-08, 1.423717e-08, 1.423203e-08, 1.423724e-08, 1.421116e-08, 
    1.422233e-08, 1.419938e-08, 1.410995e-08, 1.413624e-08, 1.405782e-08, 
    1.401064e-08, 1.397931e-08, 1.395706e-08, 1.396021e-08, 1.39662e-08, 
    1.3997e-08, 1.402596e-08, 1.404803e-08, 1.406278e-08, 1.407732e-08, 
    1.41213e-08, 1.414459e-08, 1.419671e-08, 1.418731e-08, 1.420323e-08, 
    1.421845e-08, 1.4244e-08, 1.423979e-08, 1.425104e-08, 1.420282e-08, 
    1.423487e-08, 1.418195e-08, 1.419643e-08, 1.408125e-08, 1.403738e-08, 
    1.401871e-08, 1.400238e-08, 1.396263e-08, 1.399008e-08, 1.397926e-08, 
    1.4005e-08, 1.402136e-08, 1.401327e-08, 1.406319e-08, 1.404378e-08, 
    1.414597e-08, 1.410196e-08, 1.421668e-08, 1.418924e-08, 1.422326e-08, 
    1.42059e-08, 1.423564e-08, 1.420887e-08, 1.425523e-08, 1.426532e-08, 
    1.425843e-08, 1.428492e-08, 1.420739e-08, 1.423717e-08, 1.401304e-08, 
    1.401436e-08, 1.402051e-08, 1.399348e-08, 1.399183e-08, 1.396707e-08, 
    1.398911e-08, 1.399849e-08, 1.402231e-08, 1.403639e-08, 1.404978e-08, 
    1.407921e-08, 1.411207e-08, 1.415802e-08, 1.419102e-08, 1.421313e-08, 
    1.419957e-08, 1.421154e-08, 1.419816e-08, 1.419189e-08, 1.426154e-08, 
    1.422243e-08, 1.428111e-08, 1.427787e-08, 1.425131e-08, 1.427823e-08, 
    1.401529e-08, 1.40077e-08, 1.398133e-08, 1.400196e-08, 1.396437e-08, 
    1.398541e-08, 1.399751e-08, 1.404418e-08, 1.405444e-08, 1.406394e-08, 
    1.408272e-08, 1.410681e-08, 1.414905e-08, 1.41858e-08, 1.421934e-08, 
    1.421688e-08, 1.421775e-08, 1.422524e-08, 1.420668e-08, 1.422828e-08, 
    1.423191e-08, 1.422243e-08, 1.427743e-08, 1.426172e-08, 1.42778e-08, 
    1.426757e-08, 1.401016e-08, 1.402294e-08, 1.401604e-08, 1.402901e-08, 
    1.401987e-08, 1.406052e-08, 1.407271e-08, 1.412972e-08, 1.410633e-08, 
    1.414356e-08, 1.411011e-08, 1.411604e-08, 1.414477e-08, 1.411192e-08, 
    1.418377e-08, 1.413506e-08, 1.422553e-08, 1.417689e-08, 1.422858e-08, 
    1.42192e-08, 1.423473e-08, 1.424864e-08, 1.426614e-08, 1.429841e-08, 
    1.429094e-08, 1.431793e-08, 1.404198e-08, 1.405854e-08, 1.405709e-08, 
    1.407442e-08, 1.408724e-08, 1.411502e-08, 1.415956e-08, 1.414281e-08, 
    1.417356e-08, 1.417973e-08, 1.413302e-08, 1.416169e-08, 1.406963e-08, 
    1.40845e-08, 1.407565e-08, 1.404328e-08, 1.414666e-08, 1.409362e-08, 
    1.419156e-08, 1.416284e-08, 1.424665e-08, 1.420497e-08, 1.428683e-08, 
    1.432179e-08, 1.435471e-08, 1.439315e-08, 1.406758e-08, 1.405633e-08, 
    1.407648e-08, 1.410435e-08, 1.413022e-08, 1.416459e-08, 1.416811e-08, 
    1.417454e-08, 1.419122e-08, 1.420524e-08, 1.417657e-08, 1.420875e-08, 
    1.408795e-08, 1.415127e-08, 1.405207e-08, 1.408195e-08, 1.410271e-08, 
    1.409361e-08, 1.41409e-08, 1.415204e-08, 1.419731e-08, 1.417391e-08, 
    1.431316e-08, 1.425157e-08, 1.442243e-08, 1.43747e-08, 1.40524e-08, 
    1.406755e-08, 1.412025e-08, 1.409518e-08, 1.416688e-08, 1.418453e-08, 
    1.419887e-08, 1.42172e-08, 1.421918e-08, 1.423004e-08, 1.421224e-08, 
    1.422934e-08, 1.416466e-08, 1.419357e-08, 1.411423e-08, 1.413355e-08, 
    1.412466e-08, 1.411492e-08, 1.414499e-08, 1.417702e-08, 1.417772e-08, 
    1.418798e-08, 1.42169e-08, 1.416717e-08, 1.432109e-08, 1.422605e-08, 
    1.408406e-08, 1.411323e-08, 1.41174e-08, 1.41061e-08, 1.418276e-08, 
    1.415499e-08, 1.422977e-08, 1.420957e-08, 1.424268e-08, 1.422622e-08, 
    1.42238e-08, 1.420267e-08, 1.418951e-08, 1.415626e-08, 1.41292e-08, 
    1.410774e-08, 1.411273e-08, 1.41363e-08, 1.417899e-08, 1.421936e-08, 
    1.421051e-08, 1.424016e-08, 1.416169e-08, 1.419459e-08, 1.418187e-08, 
    1.421504e-08, 1.414237e-08, 1.420423e-08, 1.412654e-08, 1.413336e-08, 
    1.415444e-08, 1.419682e-08, 1.420621e-08, 1.421621e-08, 1.421004e-08, 
    1.418007e-08, 1.417516e-08, 1.415393e-08, 1.414806e-08, 1.413188e-08, 
    1.411847e-08, 1.413072e-08, 1.414357e-08, 1.418008e-08, 1.421298e-08, 
    1.424883e-08, 1.425761e-08, 1.429947e-08, 1.426539e-08, 1.432162e-08, 
    1.42738e-08, 1.435658e-08, 1.420783e-08, 1.427241e-08, 1.41554e-08, 
    1.416801e-08, 1.419081e-08, 1.424311e-08, 1.421488e-08, 1.424789e-08, 
    1.417497e-08, 1.413711e-08, 1.412732e-08, 1.410905e-08, 1.412774e-08, 
    1.412622e-08, 1.414411e-08, 1.413836e-08, 1.41813e-08, 1.415824e-08, 
    1.422374e-08, 1.424764e-08, 1.43151e-08, 1.435644e-08, 1.439852e-08, 
    1.441709e-08, 1.442274e-08, 1.44251e-08 ;

 SOIL1N_TO_SOIL3N =
  1.657348e-10, 1.661885e-10, 1.661003e-10, 1.664662e-10, 1.662633e-10, 
    1.665028e-10, 1.658268e-10, 1.662065e-10, 1.659641e-10, 1.657757e-10, 
    1.671759e-10, 1.664825e-10, 1.678961e-10, 1.674541e-10, 1.685644e-10, 
    1.678273e-10, 1.68713e-10, 1.685432e-10, 1.690544e-10, 1.68908e-10, 
    1.695614e-10, 1.69122e-10, 1.699002e-10, 1.694565e-10, 1.695259e-10, 
    1.691075e-10, 1.666222e-10, 1.670896e-10, 1.665944e-10, 1.666611e-10, 
    1.666312e-10, 1.662675e-10, 1.660841e-10, 1.657001e-10, 1.657699e-10, 
    1.660519e-10, 1.666911e-10, 1.664742e-10, 1.670209e-10, 1.670086e-10, 
    1.676171e-10, 1.673427e-10, 1.683652e-10, 1.680747e-10, 1.689141e-10, 
    1.68703e-10, 1.689042e-10, 1.688432e-10, 1.689049e-10, 1.685954e-10, 
    1.68728e-10, 1.684556e-10, 1.673941e-10, 1.677061e-10, 1.667753e-10, 
    1.662153e-10, 1.658435e-10, 1.655795e-10, 1.656168e-10, 1.656879e-10, 
    1.660535e-10, 1.663972e-10, 1.666591e-10, 1.668343e-10, 1.670068e-10, 
    1.675289e-10, 1.678053e-10, 1.684239e-10, 1.683123e-10, 1.685013e-10, 
    1.68682e-10, 1.689852e-10, 1.689353e-10, 1.690688e-10, 1.684964e-10, 
    1.688768e-10, 1.682487e-10, 1.684206e-10, 1.670535e-10, 1.665327e-10, 
    1.663111e-10, 1.661173e-10, 1.656455e-10, 1.659713e-10, 1.658429e-10, 
    1.661484e-10, 1.663426e-10, 1.662466e-10, 1.66839e-10, 1.666087e-10, 
    1.678216e-10, 1.672993e-10, 1.686609e-10, 1.683352e-10, 1.68739e-10, 
    1.68533e-10, 1.688859e-10, 1.685683e-10, 1.691186e-10, 1.692383e-10, 
    1.691565e-10, 1.69471e-10, 1.685507e-10, 1.689041e-10, 1.662439e-10, 
    1.662595e-10, 1.663325e-10, 1.660117e-10, 1.659921e-10, 1.656982e-10, 
    1.659598e-10, 1.660711e-10, 1.663538e-10, 1.66521e-10, 1.666799e-10, 
    1.670293e-10, 1.674193e-10, 1.679646e-10, 1.683563e-10, 1.686188e-10, 
    1.684579e-10, 1.686e-10, 1.684411e-10, 1.683667e-10, 1.691935e-10, 
    1.687292e-10, 1.694258e-10, 1.693872e-10, 1.69072e-10, 1.693916e-10, 
    1.662705e-10, 1.661804e-10, 1.658675e-10, 1.661124e-10, 1.656662e-10, 
    1.659159e-10, 1.660595e-10, 1.666135e-10, 1.667352e-10, 1.66848e-10, 
    1.670709e-10, 1.673568e-10, 1.678582e-10, 1.682944e-10, 1.686925e-10, 
    1.686634e-10, 1.686736e-10, 1.687625e-10, 1.685423e-10, 1.687987e-10, 
    1.688417e-10, 1.687292e-10, 1.693821e-10, 1.691956e-10, 1.693864e-10, 
    1.69265e-10, 1.662097e-10, 1.663613e-10, 1.662794e-10, 1.664335e-10, 
    1.663249e-10, 1.668074e-10, 1.669521e-10, 1.676288e-10, 1.673511e-10, 
    1.67793e-10, 1.67396e-10, 1.674664e-10, 1.678074e-10, 1.674175e-10, 
    1.682703e-10, 1.676921e-10, 1.68766e-10, 1.681887e-10, 1.688022e-10, 
    1.686908e-10, 1.688752e-10, 1.690403e-10, 1.69248e-10, 1.696311e-10, 
    1.695424e-10, 1.698628e-10, 1.665874e-10, 1.667839e-10, 1.667667e-10, 
    1.669724e-10, 1.671245e-10, 1.674542e-10, 1.679829e-10, 1.677841e-10, 
    1.681491e-10, 1.682223e-10, 1.676679e-10, 1.680083e-10, 1.669155e-10, 
    1.670921e-10, 1.66987e-10, 1.666028e-10, 1.678299e-10, 1.672002e-10, 
    1.683628e-10, 1.680218e-10, 1.690167e-10, 1.68522e-10, 1.694936e-10, 
    1.699086e-10, 1.702994e-10, 1.707557e-10, 1.668913e-10, 1.667577e-10, 
    1.669969e-10, 1.673277e-10, 1.676347e-10, 1.680426e-10, 1.680844e-10, 
    1.681608e-10, 1.683587e-10, 1.685251e-10, 1.681849e-10, 1.685668e-10, 
    1.671329e-10, 1.678845e-10, 1.667071e-10, 1.670617e-10, 1.673082e-10, 
    1.672001e-10, 1.677614e-10, 1.678937e-10, 1.68431e-10, 1.681533e-10, 
    1.698062e-10, 1.690751e-10, 1.711032e-10, 1.705366e-10, 1.66711e-10, 
    1.668908e-10, 1.675164e-10, 1.672188e-10, 1.680699e-10, 1.682793e-10, 
    1.684495e-10, 1.686671e-10, 1.686906e-10, 1.688195e-10, 1.686083e-10, 
    1.688112e-10, 1.680435e-10, 1.683866e-10, 1.674449e-10, 1.676742e-10, 
    1.675687e-10, 1.674531e-10, 1.678101e-10, 1.681902e-10, 1.681984e-10, 
    1.683203e-10, 1.686636e-10, 1.680733e-10, 1.699003e-10, 1.687721e-10, 
    1.670869e-10, 1.67433e-10, 1.674825e-10, 1.673484e-10, 1.682583e-10, 
    1.679287e-10, 1.688164e-10, 1.685765e-10, 1.689695e-10, 1.687742e-10, 
    1.687455e-10, 1.684947e-10, 1.683385e-10, 1.679438e-10, 1.676226e-10, 
    1.673679e-10, 1.674271e-10, 1.677069e-10, 1.682135e-10, 1.686927e-10, 
    1.685877e-10, 1.689396e-10, 1.680082e-10, 1.683988e-10, 1.682478e-10, 
    1.686415e-10, 1.677789e-10, 1.685132e-10, 1.675911e-10, 1.676719e-10, 
    1.679221e-10, 1.684252e-10, 1.685366e-10, 1.686554e-10, 1.685821e-10, 
    1.682264e-10, 1.681681e-10, 1.679161e-10, 1.678464e-10, 1.676543e-10, 
    1.674953e-10, 1.676406e-10, 1.677932e-10, 1.682266e-10, 1.68617e-10, 
    1.690426e-10, 1.691468e-10, 1.696437e-10, 1.692391e-10, 1.699066e-10, 
    1.69339e-10, 1.703216e-10, 1.685559e-10, 1.693224e-10, 1.679335e-10, 
    1.680832e-10, 1.683539e-10, 1.689746e-10, 1.686396e-10, 1.690314e-10, 
    1.681659e-10, 1.677165e-10, 1.676003e-10, 1.673834e-10, 1.676053e-10, 
    1.675872e-10, 1.677996e-10, 1.677313e-10, 1.68241e-10, 1.679672e-10, 
    1.687448e-10, 1.690284e-10, 1.698292e-10, 1.703199e-10, 1.708194e-10, 
    1.710398e-10, 1.711069e-10, 1.711349e-10 ;

 SOIL1N_vr =
  2.497551, 2.497545, 2.497546, 2.497541, 2.497544, 2.497541, 2.49755, 
    2.497545, 2.497548, 2.497551, 2.497531, 2.497541, 2.497521, 2.497528, 
    2.497512, 2.497522, 2.49751, 2.497513, 2.497505, 2.497507, 2.497499, 
    2.497504, 2.497494, 2.4975, 2.497499, 2.497505, 2.497539, 2.497533, 
    2.497539, 2.497539, 2.497539, 2.497544, 2.497546, 2.497552, 2.497551, 
    2.497547, 2.497538, 2.497541, 2.497534, 2.497534, 2.497525, 2.497529, 
    2.497515, 2.497519, 2.497507, 2.49751, 2.497508, 2.497508, 2.497508, 
    2.497512, 2.49751, 2.497514, 2.497528, 2.497524, 2.497537, 2.497545, 
    2.49755, 2.497553, 2.497553, 2.497552, 2.497547, 2.497542, 2.497539, 
    2.497536, 2.497534, 2.497526, 2.497523, 2.497514, 2.497516, 2.497513, 
    2.49751, 2.497506, 2.497507, 2.497505, 2.497513, 2.497508, 2.497517, 
    2.497514, 2.497533, 2.49754, 2.497543, 2.497546, 2.497553, 2.497548, 
    2.49755, 2.497545, 2.497543, 2.497544, 2.497536, 2.497539, 2.497522, 
    2.49753, 2.497511, 2.497515, 2.49751, 2.497513, 2.497508, 2.497512, 
    2.497504, 2.497503, 2.497504, 2.4975, 2.497512, 2.497508, 2.497544, 
    2.497544, 2.497543, 2.497547, 2.497548, 2.497552, 2.497548, 2.497547, 
    2.497543, 2.49754, 2.497538, 2.497533, 2.497528, 2.49752, 2.497515, 
    2.497511, 2.497514, 2.497512, 2.497514, 2.497515, 2.497504, 2.49751, 
    2.4975, 2.497501, 2.497505, 2.497501, 2.497544, 2.497545, 2.49755, 
    2.497546, 2.497552, 2.497549, 2.497547, 2.497539, 2.497537, 2.497536, 
    2.497533, 2.497529, 2.497522, 2.497516, 2.49751, 2.497511, 2.497511, 
    2.497509, 2.497513, 2.497509, 2.497508, 2.49751, 2.497501, 2.497504, 
    2.497501, 2.497503, 2.497545, 2.497543, 2.497544, 2.497542, 2.497543, 
    2.497536, 2.497535, 2.497525, 2.497529, 2.497523, 2.497528, 2.497527, 
    2.497523, 2.497528, 2.497516, 2.497524, 2.497509, 2.497517, 2.497509, 
    2.49751, 2.497508, 2.497506, 2.497503, 2.497498, 2.497499, 2.497494, 
    2.49754, 2.497537, 2.497537, 2.497534, 2.497532, 2.497528, 2.49752, 
    2.497523, 2.497518, 2.497517, 2.497524, 2.49752, 2.497535, 2.497533, 
    2.497534, 2.497539, 2.497522, 2.497531, 2.497515, 2.49752, 2.497506, 
    2.497513, 2.497499, 2.497494, 2.497488, 2.497482, 2.497535, 2.497537, 
    2.497534, 2.497529, 2.497525, 2.497519, 2.497519, 2.497518, 2.497515, 
    2.497513, 2.497517, 2.497512, 2.497532, 2.497522, 2.497538, 2.497533, 
    2.49753, 2.497531, 2.497523, 2.497521, 2.497514, 2.497518, 2.497495, 
    2.497505, 2.497477, 2.497485, 2.497538, 2.497535, 2.497527, 2.497531, 
    2.497519, 2.497516, 2.497514, 2.497511, 2.49751, 2.497509, 2.497512, 
    2.497509, 2.497519, 2.497515, 2.497528, 2.497524, 2.497526, 2.497528, 
    2.497523, 2.497517, 2.497517, 2.497515, 2.497511, 2.497519, 2.497494, 
    2.497509, 2.497533, 2.497528, 2.497527, 2.497529, 2.497516, 2.497521, 
    2.497509, 2.497512, 2.497507, 2.497509, 2.49751, 2.497513, 2.497515, 
    2.497521, 2.497525, 2.497529, 2.497528, 2.497524, 2.497517, 2.49751, 
    2.497512, 2.497507, 2.49752, 2.497514, 2.497517, 2.497511, 2.497523, 
    2.497513, 2.497526, 2.497524, 2.497521, 2.497514, 2.497513, 2.497511, 
    2.497512, 2.497517, 2.497518, 2.497521, 2.497522, 2.497525, 2.497527, 
    2.497525, 2.497523, 2.497517, 2.497511, 2.497506, 2.497504, 2.497497, 
    2.497503, 2.497494, 2.497502, 2.497488, 2.497512, 2.497502, 2.497521, 
    2.497519, 2.497515, 2.497507, 2.497511, 2.497506, 2.497518, 2.497524, 
    2.497525, 2.497529, 2.497525, 2.497526, 2.497523, 2.497524, 2.497517, 
    2.49752, 2.49751, 2.497506, 2.497495, 2.497488, 2.497481, 2.497478, 
    2.497477, 2.497477,
  2.497528, 2.497521, 2.497523, 2.497517, 2.49752, 2.497517, 2.497527, 
    2.497521, 2.497525, 2.497527, 2.497507, 2.497517, 2.497497, 2.497503, 
    2.497487, 2.497498, 2.497485, 2.497488, 2.49748, 2.497483, 2.497473, 
    2.497479, 2.497468, 2.497475, 2.497473, 2.49748, 2.497515, 2.497509, 
    2.497516, 2.497515, 2.497515, 2.49752, 2.497523, 2.497528, 2.497527, 
    2.497523, 2.497514, 2.497517, 2.497509, 2.49751, 2.497501, 2.497505, 
    2.49749, 2.497494, 2.497482, 2.497485, 2.497483, 2.497483, 2.497483, 
    2.497487, 2.497485, 2.497489, 2.497504, 2.4975, 2.497513, 2.497521, 
    2.497526, 2.49753, 2.49753, 2.497529, 2.497523, 2.497518, 2.497515, 
    2.497512, 2.49751, 2.497502, 2.497498, 2.497489, 2.497491, 2.497488, 
    2.497486, 2.497481, 2.497482, 2.49748, 2.497488, 2.497483, 2.497492, 
    2.497489, 2.497509, 2.497516, 2.49752, 2.497522, 2.497529, 2.497524, 
    2.497526, 2.497522, 2.497519, 2.497521, 2.497512, 2.497515, 2.497498, 
    2.497505, 2.497486, 2.497491, 2.497485, 2.497488, 2.497483, 2.497487, 
    2.497479, 2.497478, 2.497479, 2.497474, 2.497488, 2.497483, 2.497521, 
    2.49752, 2.497519, 2.497524, 2.497524, 2.497529, 2.497525, 2.497523, 
    2.497519, 2.497517, 2.497514, 2.497509, 2.497504, 2.497496, 2.49749, 
    2.497487, 2.497489, 2.497487, 2.497489, 2.49749, 2.497478, 2.497485, 
    2.497475, 2.497476, 2.49748, 2.497476, 2.49752, 2.497522, 2.497526, 
    2.497523, 2.497529, 2.497525, 2.497523, 2.497515, 2.497514, 2.497512, 
    2.497509, 2.497505, 2.497498, 2.497491, 2.497485, 2.497486, 2.497486, 
    2.497484, 2.497488, 2.497484, 2.497483, 2.497485, 2.497476, 2.497478, 
    2.497476, 2.497477, 2.497521, 2.497519, 2.49752, 2.497518, 2.497519, 
    2.497513, 2.49751, 2.497501, 2.497505, 2.497498, 2.497504, 2.497503, 
    2.497498, 2.497504, 2.497492, 2.4975, 2.497484, 2.497493, 2.497484, 
    2.497486, 2.497483, 2.497481, 2.497478, 2.497472, 2.497473, 2.497469, 
    2.497516, 2.497513, 2.497513, 2.49751, 2.497508, 2.497503, 2.497496, 
    2.497499, 2.497493, 2.497492, 2.4975, 2.497495, 2.497511, 2.497509, 
    2.49751, 2.497515, 2.497498, 2.497507, 2.49749, 2.497495, 2.497481, 
    2.497488, 2.497474, 2.497468, 2.497463, 2.497456, 2.497511, 2.497513, 
    2.49751, 2.497505, 2.497501, 2.497495, 2.497494, 2.497493, 2.49749, 
    2.497488, 2.497493, 2.497487, 2.497508, 2.497497, 2.497514, 2.497509, 
    2.497505, 2.497507, 2.497499, 2.497497, 2.497489, 2.497493, 2.49747, 
    2.49748, 2.497451, 2.497459, 2.497514, 2.497511, 2.497502, 2.497507, 
    2.497494, 2.497491, 2.497489, 2.497486, 2.497486, 2.497484, 2.497487, 
    2.497484, 2.497495, 2.49749, 2.497503, 2.4975, 2.497502, 2.497503, 
    2.497498, 2.497493, 2.497493, 2.497491, 2.497486, 2.497494, 2.497468, 
    2.497484, 2.497509, 2.497504, 2.497503, 2.497505, 2.497492, 2.497496, 
    2.497484, 2.497487, 2.497482, 2.497484, 2.497485, 2.497488, 2.497491, 
    2.497496, 2.497501, 2.497504, 2.497504, 2.4975, 2.497492, 2.497485, 
    2.497487, 2.497482, 2.497495, 2.49749, 2.497492, 2.497486, 2.497499, 
    2.497488, 2.497501, 2.4975, 2.497497, 2.497489, 2.497488, 2.497486, 
    2.497487, 2.497492, 2.497493, 2.497497, 2.497498, 2.4975, 2.497503, 
    2.497501, 2.497498, 2.497492, 2.497487, 2.49748, 2.497479, 2.497472, 
    2.497478, 2.497468, 2.497476, 2.497462, 2.497488, 2.497477, 2.497496, 
    2.497494, 2.49749, 2.497482, 2.497486, 2.497481, 2.497493, 2.497499, 
    2.497501, 2.497504, 2.497501, 2.497501, 2.497498, 2.497499, 2.497492, 
    2.497496, 2.497485, 2.497481, 2.497469, 2.497462, 2.497455, 2.497452, 
    2.497451, 2.497451,
  2.49752, 2.497513, 2.497514, 2.497509, 2.497512, 2.497509, 2.497519, 
    2.497513, 2.497516, 2.497519, 2.497499, 2.497509, 2.497488, 2.497495, 
    2.497479, 2.497489, 2.497477, 2.497479, 2.497472, 2.497474, 2.497464, 
    2.497471, 2.497459, 2.497466, 2.497465, 2.497471, 2.497507, 2.4975, 
    2.497507, 2.497506, 2.497507, 2.497512, 2.497515, 2.49752, 2.497519, 
    2.497515, 2.497506, 2.497509, 2.497501, 2.497501, 2.497492, 2.497496, 
    2.497482, 2.497486, 2.497473, 2.497477, 2.497474, 2.497475, 2.497474, 
    2.497478, 2.497476, 2.49748, 2.497496, 2.497491, 2.497505, 2.497513, 
    2.497518, 2.497522, 2.497522, 2.49752, 2.497515, 2.49751, 2.497506, 
    2.497504, 2.497501, 2.497494, 2.49749, 2.497481, 2.497482, 2.49748, 
    2.497477, 2.497473, 2.497473, 2.497471, 2.49748, 2.497474, 2.497483, 
    2.497481, 2.497501, 2.497508, 2.497511, 2.497514, 2.497521, 2.497516, 
    2.497518, 2.497514, 2.497511, 2.497512, 2.497504, 2.497507, 2.497489, 
    2.497497, 2.497477, 2.497482, 2.497476, 2.497479, 2.497474, 2.497479, 
    2.497471, 2.497469, 2.49747, 2.497466, 2.497479, 2.497474, 2.497512, 
    2.497512, 2.497511, 2.497516, 2.497516, 2.49752, 2.497517, 2.497515, 
    2.497511, 2.497508, 2.497506, 2.497501, 2.497495, 2.497487, 2.497482, 
    2.497478, 2.49748, 2.497478, 2.49748, 2.497482, 2.497469, 2.497476, 
    2.497466, 2.497467, 2.497471, 2.497467, 2.497512, 2.497513, 2.497518, 
    2.497514, 2.497521, 2.497517, 2.497515, 2.497507, 2.497505, 2.497504, 
    2.4975, 2.497496, 2.497489, 2.497483, 2.497477, 2.497477, 2.497477, 
    2.497476, 2.497479, 2.497475, 2.497475, 2.497476, 2.497467, 2.497469, 
    2.497467, 2.497468, 2.497513, 2.497511, 2.497512, 2.49751, 2.497511, 
    2.497504, 2.497502, 2.497492, 2.497496, 2.49749, 2.497496, 2.497495, 
    2.49749, 2.497495, 2.497483, 2.497491, 2.497476, 2.497484, 2.497475, 
    2.497477, 2.497474, 2.497472, 2.497469, 2.497463, 2.497464, 2.49746, 
    2.497507, 2.497504, 2.497505, 2.497502, 2.4975, 2.497495, 2.497487, 
    2.49749, 2.497485, 2.497484, 2.497492, 2.497487, 2.497503, 2.4975, 
    2.497502, 2.497507, 2.497489, 2.497499, 2.497482, 2.497487, 2.497472, 
    2.497479, 2.497465, 2.497459, 2.497453, 2.497447, 2.497503, 2.497505, 
    2.497501, 2.497497, 2.497492, 2.497486, 2.497486, 2.497484, 2.497482, 
    2.497479, 2.497484, 2.497479, 2.497499, 2.497488, 2.497506, 2.4975, 
    2.497497, 2.497499, 2.49749, 2.497488, 2.497481, 2.497485, 2.497461, 
    2.497471, 2.497442, 2.49745, 2.497506, 2.497503, 2.497494, 2.497498, 
    2.497486, 2.497483, 2.49748, 2.497477, 2.497477, 2.497475, 2.497478, 
    2.497475, 2.497486, 2.497481, 2.497495, 2.497492, 2.497493, 2.497495, 
    2.49749, 2.497484, 2.497484, 2.497482, 2.497477, 2.497486, 2.497459, 
    2.497476, 2.4975, 2.497495, 2.497494, 2.497496, 2.497483, 2.497488, 
    2.497475, 2.497478, 2.497473, 2.497476, 2.497476, 2.49748, 2.497482, 
    2.497488, 2.497492, 2.497496, 2.497495, 2.497491, 2.497484, 2.497477, 
    2.497478, 2.497473, 2.497487, 2.497481, 2.497483, 2.497478, 2.49749, 
    2.497479, 2.497493, 2.497492, 2.497488, 2.497481, 2.497479, 2.497477, 
    2.497478, 2.497483, 2.497484, 2.497488, 2.497489, 2.497492, 2.497494, 
    2.497492, 2.49749, 2.497483, 2.497478, 2.497472, 2.49747, 2.497463, 
    2.497469, 2.497459, 2.497468, 2.497453, 2.497479, 2.497468, 2.497488, 
    2.497486, 2.497482, 2.497473, 2.497478, 2.497472, 2.497484, 2.497491, 
    2.497493, 2.497496, 2.497493, 2.497493, 2.49749, 2.497491, 2.497483, 
    2.497487, 2.497476, 2.497472, 2.49746, 2.497453, 2.497446, 2.497443, 
    2.497442, 2.497442,
  2.497596, 2.497589, 2.49759, 2.497585, 2.497588, 2.497585, 2.497594, 
    2.497589, 2.497592, 2.497595, 2.497575, 2.497585, 2.497565, 2.497571, 
    2.497555, 2.497566, 2.497553, 2.497555, 2.497548, 2.49755, 2.497541, 
    2.497547, 2.497536, 2.497542, 2.497541, 2.497547, 2.497583, 2.497576, 
    2.497583, 2.497582, 2.497583, 2.497588, 2.497591, 2.497596, 2.497595, 
    2.497591, 2.497582, 2.497585, 2.497577, 2.497577, 2.497569, 2.497572, 
    2.497558, 2.497562, 2.49755, 2.497553, 2.49755, 2.497551, 2.49755, 
    2.497555, 2.497553, 2.497556, 2.497572, 2.497567, 2.497581, 2.497589, 
    2.497594, 2.497598, 2.497597, 2.497596, 2.497591, 2.497586, 2.497582, 
    2.49758, 2.497577, 2.49757, 2.497566, 2.497557, 2.497559, 2.497556, 
    2.497553, 2.497549, 2.49755, 2.497548, 2.497556, 2.49755, 2.49756, 
    2.497557, 2.497577, 2.497584, 2.497587, 2.49759, 2.497597, 2.497592, 
    2.497594, 2.49759, 2.497587, 2.497588, 2.49758, 2.497583, 2.497566, 
    2.497573, 2.497554, 2.497558, 2.497552, 2.497555, 2.49755, 2.497555, 
    2.497547, 2.497545, 2.497546, 2.497542, 2.497555, 2.49755, 2.497588, 
    2.497588, 2.497587, 2.497591, 2.497592, 2.497596, 2.497592, 2.497591, 
    2.497587, 2.497584, 2.497582, 2.497577, 2.497571, 2.497564, 2.497558, 
    2.497554, 2.497556, 2.497554, 2.497557, 2.497558, 2.497546, 2.497553, 
    2.497543, 2.497543, 2.497548, 2.497543, 2.497588, 2.497589, 2.497594, 
    2.49759, 2.497597, 2.497593, 2.497591, 2.497583, 2.497581, 2.49758, 
    2.497576, 2.497572, 2.497565, 2.497559, 2.497553, 2.497554, 2.497553, 
    2.497552, 2.497555, 2.497552, 2.497551, 2.497553, 2.497543, 2.497546, 
    2.497543, 2.497545, 2.497589, 2.497586, 2.497588, 2.497586, 2.497587, 
    2.49758, 2.497578, 2.497568, 2.497572, 2.497566, 2.497572, 2.497571, 
    2.497566, 2.497571, 2.497559, 2.497567, 2.497552, 2.49756, 2.497551, 
    2.497553, 2.49755, 2.497548, 2.497545, 2.49754, 2.497541, 2.497536, 
    2.497583, 2.497581, 2.497581, 2.497578, 2.497576, 2.497571, 2.497563, 
    2.497566, 2.497561, 2.49756, 2.497568, 2.497563, 2.497579, 2.497576, 
    2.497578, 2.497583, 2.497566, 2.497575, 2.497558, 2.497563, 2.497548, 
    2.497555, 2.497542, 2.497536, 2.49753, 2.497524, 2.497579, 2.497581, 
    2.497577, 2.497573, 2.497568, 2.497562, 2.497562, 2.497561, 2.497558, 
    2.497555, 2.49756, 2.497555, 2.497576, 2.497565, 2.497582, 2.497576, 
    2.497573, 2.497575, 2.497566, 2.497565, 2.497557, 2.497561, 2.497537, 
    2.497548, 2.497519, 2.497527, 2.497581, 2.497579, 2.49757, 2.497574, 
    2.497562, 2.497559, 2.497557, 2.497553, 2.497553, 2.497551, 2.497554, 
    2.497551, 2.497562, 2.497557, 2.497571, 2.497568, 2.497569, 2.497571, 
    2.497566, 2.49756, 2.49756, 2.497558, 2.497554, 2.497562, 2.497536, 
    2.497552, 2.497576, 2.497571, 2.497571, 2.497572, 2.497559, 2.497564, 
    2.497551, 2.497555, 2.497549, 2.497552, 2.497552, 2.497556, 2.497558, 
    2.497564, 2.497568, 2.497572, 2.497571, 2.497567, 2.49756, 2.497553, 
    2.497555, 2.49755, 2.497563, 2.497557, 2.49756, 2.497554, 2.497566, 
    2.497556, 2.497569, 2.497568, 2.497564, 2.497557, 2.497555, 2.497554, 
    2.497555, 2.49756, 2.497561, 2.497564, 2.497565, 2.497568, 2.49757, 
    2.497568, 2.497566, 2.49756, 2.497554, 2.497548, 2.497547, 2.49754, 
    2.497545, 2.497536, 2.497544, 2.49753, 2.497555, 2.497544, 2.497564, 
    2.497562, 2.497558, 2.497549, 2.497554, 2.497548, 2.497561, 2.497567, 
    2.497569, 2.497572, 2.497569, 2.497569, 2.497566, 2.497567, 2.49756, 
    2.497564, 2.497552, 2.497548, 2.497537, 2.49753, 2.497523, 2.497519, 
    2.497519, 2.497518,
  2.497849, 2.497843, 2.497844, 2.497839, 2.497842, 2.497839, 2.497848, 
    2.497843, 2.497846, 2.497849, 2.49783, 2.497839, 2.49782, 2.497826, 
    2.497812, 2.497821, 2.497809, 2.497812, 2.497805, 2.497807, 2.497798, 
    2.497804, 2.497793, 2.497799, 2.497799, 2.497804, 2.497837, 2.497831, 
    2.497838, 2.497837, 2.497837, 2.497842, 2.497844, 2.49785, 2.497849, 
    2.497845, 2.497837, 2.497839, 2.497832, 2.497832, 2.497824, 2.497828, 
    2.497814, 2.497818, 2.497807, 2.49781, 2.497807, 2.497808, 2.497807, 
    2.497811, 2.497809, 2.497813, 2.497827, 2.497823, 2.497835, 2.497843, 
    2.497848, 2.497851, 2.497851, 2.49785, 2.497845, 2.49784, 2.497837, 
    2.497834, 2.497832, 2.497825, 2.497822, 2.497813, 2.497815, 2.497812, 
    2.49781, 2.497806, 2.497807, 2.497805, 2.497812, 2.497807, 2.497816, 
    2.497813, 2.497832, 2.497838, 2.497842, 2.497844, 2.49785, 2.497846, 
    2.497848, 2.497844, 2.497841, 2.497842, 2.497834, 2.497838, 2.497821, 
    2.497828, 2.49781, 2.497814, 2.497809, 2.497812, 2.497807, 2.497811, 
    2.497804, 2.497802, 2.497803, 2.497799, 2.497812, 2.497807, 2.497843, 
    2.497842, 2.497841, 2.497846, 2.497846, 2.49785, 2.497846, 2.497845, 
    2.497841, 2.497839, 2.497837, 2.497832, 2.497827, 2.497819, 2.497814, 
    2.497811, 2.497813, 2.497811, 2.497813, 2.497814, 2.497803, 2.497809, 
    2.4978, 2.4978, 2.497805, 2.4978, 2.497842, 2.497843, 2.497848, 2.497844, 
    2.49785, 2.497847, 2.497845, 2.497838, 2.497836, 2.497834, 2.497831, 
    2.497828, 2.497821, 2.497815, 2.49781, 2.49781, 2.49781, 2.497809, 
    2.497812, 2.497808, 2.497808, 2.497809, 2.497801, 2.497803, 2.4978, 
    2.497802, 2.497843, 2.497841, 2.497842, 2.49784, 2.497841, 2.497835, 
    2.497833, 2.497824, 2.497828, 2.497822, 2.497827, 2.497826, 2.497822, 
    2.497827, 2.497815, 2.497823, 2.497809, 2.497817, 2.497808, 2.49781, 
    2.497807, 2.497805, 2.497802, 2.497797, 2.497798, 2.497794, 2.497838, 
    2.497835, 2.497835, 2.497833, 2.497831, 2.497826, 2.497819, 2.497822, 
    2.497817, 2.497816, 2.497823, 2.497819, 2.497833, 2.497831, 2.497833, 
    2.497838, 2.497821, 2.49783, 2.497814, 2.497819, 2.497805, 2.497812, 
    2.497799, 2.497793, 2.497788, 2.497782, 2.497834, 2.497836, 2.497832, 
    2.497828, 2.497824, 2.497818, 2.497818, 2.497817, 2.497814, 2.497812, 
    2.497817, 2.497811, 2.497831, 2.497821, 2.497836, 2.497832, 2.497828, 
    2.49783, 2.497822, 2.49782, 2.497813, 2.497817, 2.497795, 2.497805, 
    2.497777, 2.497785, 2.497836, 2.497834, 2.497825, 2.497829, 2.497818, 
    2.497815, 2.497813, 2.49781, 2.49781, 2.497808, 2.497811, 2.497808, 
    2.497818, 2.497814, 2.497826, 2.497823, 2.497825, 2.497826, 2.497822, 
    2.497817, 2.497816, 2.497815, 2.49781, 2.497818, 2.497793, 2.497809, 
    2.497831, 2.497827, 2.497826, 2.497828, 2.497816, 2.49782, 2.497808, 
    2.497811, 2.497806, 2.497809, 2.497809, 2.497812, 2.497814, 2.49782, 
    2.497824, 2.497828, 2.497827, 2.497823, 2.497816, 2.49781, 2.497811, 
    2.497806, 2.497819, 2.497814, 2.497816, 2.49781, 2.497822, 2.497812, 
    2.497824, 2.497823, 2.49782, 2.497813, 2.497812, 2.49781, 2.497811, 
    2.497816, 2.497817, 2.49782, 2.497821, 2.497824, 2.497826, 2.497824, 
    2.497822, 2.497816, 2.497811, 2.497805, 2.497804, 2.497797, 2.497802, 
    2.497793, 2.497801, 2.497788, 2.497812, 2.497801, 2.49782, 2.497818, 
    2.497814, 2.497806, 2.49781, 2.497805, 2.497817, 2.497823, 2.497824, 
    2.497827, 2.497824, 2.497824, 2.497822, 2.497823, 2.497816, 2.497819, 
    2.497809, 2.497805, 2.497794, 2.497788, 2.497781, 2.497778, 2.497777, 
    2.497777,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  7.361761e-08, 7.381911e-08, 7.377995e-08, 7.394242e-08, 7.385231e-08, 
    7.395868e-08, 7.365848e-08, 7.38271e-08, 7.371947e-08, 7.363577e-08, 
    7.425758e-08, 7.394968e-08, 7.457744e-08, 7.438113e-08, 7.48742e-08, 
    7.454688e-08, 7.494019e-08, 7.486479e-08, 7.509178e-08, 7.502676e-08, 
    7.531695e-08, 7.512179e-08, 7.546738e-08, 7.527036e-08, 7.530117e-08, 
    7.511535e-08, 7.401168e-08, 7.421925e-08, 7.399937e-08, 7.402898e-08, 
    7.40157e-08, 7.385416e-08, 7.377272e-08, 7.360223e-08, 7.363319e-08, 
    7.375842e-08, 7.404229e-08, 7.394596e-08, 7.418877e-08, 7.418329e-08, 
    7.44535e-08, 7.433168e-08, 7.478572e-08, 7.465671e-08, 7.502948e-08, 
    7.493574e-08, 7.502506e-08, 7.499798e-08, 7.502542e-08, 7.488795e-08, 
    7.494685e-08, 7.482588e-08, 7.435449e-08, 7.449304e-08, 7.407971e-08, 
    7.383102e-08, 7.366587e-08, 7.354863e-08, 7.356521e-08, 7.35968e-08, 
    7.375915e-08, 7.39118e-08, 7.402809e-08, 7.410587e-08, 7.41825e-08, 
    7.441433e-08, 7.453708e-08, 7.481178e-08, 7.476225e-08, 7.484619e-08, 
    7.492642e-08, 7.506105e-08, 7.50389e-08, 7.50982e-08, 7.4844e-08, 
    7.501294e-08, 7.473402e-08, 7.481031e-08, 7.420323e-08, 7.397196e-08, 
    7.387354e-08, 7.378748e-08, 7.357795e-08, 7.372264e-08, 7.36656e-08, 
    7.380132e-08, 7.388752e-08, 7.384489e-08, 7.410799e-08, 7.400572e-08, 
    7.454435e-08, 7.431239e-08, 7.491705e-08, 7.477242e-08, 7.495173e-08, 
    7.486024e-08, 7.501698e-08, 7.487592e-08, 7.512028e-08, 7.517347e-08, 
    7.513712e-08, 7.527677e-08, 7.48681e-08, 7.502506e-08, 7.384369e-08, 
    7.385064e-08, 7.388304e-08, 7.374061e-08, 7.37319e-08, 7.360138e-08, 
    7.371753e-08, 7.376698e-08, 7.389253e-08, 7.396677e-08, 7.403733e-08, 
    7.419247e-08, 7.436568e-08, 7.460784e-08, 7.478179e-08, 7.489836e-08, 
    7.482689e-08, 7.488999e-08, 7.481945e-08, 7.478639e-08, 7.515353e-08, 
    7.494739e-08, 7.525669e-08, 7.523958e-08, 7.509961e-08, 7.524151e-08, 
    7.385553e-08, 7.381552e-08, 7.367655e-08, 7.378531e-08, 7.358716e-08, 
    7.369807e-08, 7.376183e-08, 7.400783e-08, 7.406189e-08, 7.411199e-08, 
    7.421095e-08, 7.433791e-08, 7.456059e-08, 7.475428e-08, 7.493109e-08, 
    7.491813e-08, 7.49227e-08, 7.496217e-08, 7.486437e-08, 7.497823e-08, 
    7.499733e-08, 7.494738e-08, 7.523729e-08, 7.515448e-08, 7.523922e-08, 
    7.518531e-08, 7.382853e-08, 7.389585e-08, 7.385947e-08, 7.392788e-08, 
    7.387968e-08, 7.409395e-08, 7.415819e-08, 7.44587e-08, 7.433541e-08, 
    7.453165e-08, 7.435536e-08, 7.438658e-08, 7.4538e-08, 7.436489e-08, 
    7.474358e-08, 7.448683e-08, 7.496371e-08, 7.470734e-08, 7.497977e-08, 
    7.493033e-08, 7.50122e-08, 7.508551e-08, 7.517775e-08, 7.534788e-08, 
    7.53085e-08, 7.545077e-08, 7.399623e-08, 7.408352e-08, 7.407586e-08, 
    7.416721e-08, 7.423477e-08, 7.43812e-08, 7.461596e-08, 7.45277e-08, 
    7.468976e-08, 7.472228e-08, 7.447608e-08, 7.462723e-08, 7.414196e-08, 
    7.422036e-08, 7.417369e-08, 7.40031e-08, 7.454801e-08, 7.42684e-08, 
    7.478466e-08, 7.463326e-08, 7.507506e-08, 7.485535e-08, 7.528681e-08, 
    7.547112e-08, 7.564465e-08, 7.584727e-08, 7.413118e-08, 7.407187e-08, 
    7.417809e-08, 7.432498e-08, 7.446131e-08, 7.464248e-08, 7.466103e-08, 
    7.469496e-08, 7.478286e-08, 7.485675e-08, 7.470567e-08, 7.487527e-08, 
    7.423851e-08, 7.457228e-08, 7.404942e-08, 7.420688e-08, 7.431633e-08, 
    7.426834e-08, 7.451762e-08, 7.457635e-08, 7.481496e-08, 7.469163e-08, 
    7.542562e-08, 7.510097e-08, 7.600158e-08, 7.574999e-08, 7.405114e-08, 
    7.413099e-08, 7.440879e-08, 7.427663e-08, 7.465459e-08, 7.474758e-08, 
    7.482319e-08, 7.49198e-08, 7.493024e-08, 7.498747e-08, 7.489368e-08, 
    7.498377e-08, 7.464287e-08, 7.479523e-08, 7.437707e-08, 7.447886e-08, 
    7.443204e-08, 7.438067e-08, 7.453921e-08, 7.470804e-08, 7.471168e-08, 
    7.47658e-08, 7.491823e-08, 7.465612e-08, 7.546745e-08, 7.496644e-08, 
    7.421805e-08, 7.437176e-08, 7.439375e-08, 7.433421e-08, 7.473826e-08, 
    7.459188e-08, 7.498608e-08, 7.487957e-08, 7.505409e-08, 7.496737e-08, 
    7.495461e-08, 7.484322e-08, 7.477385e-08, 7.459859e-08, 7.445595e-08, 
    7.434285e-08, 7.436915e-08, 7.449339e-08, 7.471838e-08, 7.493117e-08, 
    7.488456e-08, 7.504082e-08, 7.462719e-08, 7.480065e-08, 7.47336e-08, 
    7.490841e-08, 7.452535e-08, 7.485146e-08, 7.444195e-08, 7.447787e-08, 
    7.458897e-08, 7.481238e-08, 7.486186e-08, 7.491461e-08, 7.488207e-08, 
    7.472409e-08, 7.469822e-08, 7.458628e-08, 7.455535e-08, 7.447006e-08, 
    7.439941e-08, 7.446395e-08, 7.453171e-08, 7.472417e-08, 7.489756e-08, 
    7.508655e-08, 7.513281e-08, 7.535348e-08, 7.517381e-08, 7.547023e-08, 
    7.521816e-08, 7.56545e-08, 7.487041e-08, 7.52108e-08, 7.459404e-08, 
    7.466052e-08, 7.478071e-08, 7.505636e-08, 7.49076e-08, 7.508159e-08, 
    7.46972e-08, 7.449766e-08, 7.444606e-08, 7.434972e-08, 7.444827e-08, 
    7.444025e-08, 7.453454e-08, 7.450424e-08, 7.473056e-08, 7.460901e-08, 
    7.495428e-08, 7.508023e-08, 7.543585e-08, 7.565375e-08, 7.587555e-08, 
    7.597343e-08, 7.600323e-08, 7.601568e-08 ;

 SOIL1_HR_S3 =
  8.7353e-10, 8.75922e-10, 8.754572e-10, 8.773859e-10, 8.763162e-10, 
    8.77579e-10, 8.740151e-10, 8.760168e-10, 8.747392e-10, 8.737456e-10, 
    8.811274e-10, 8.774721e-10, 8.849246e-10, 8.825941e-10, 8.884478e-10, 
    8.845619e-10, 8.892312e-10, 8.883361e-10, 8.910309e-10, 8.90259e-10, 
    8.937041e-10, 8.913871e-10, 8.954901e-10, 8.931511e-10, 8.935169e-10, 
    8.913106e-10, 8.782082e-10, 8.806723e-10, 8.78062e-10, 8.784135e-10, 
    8.782559e-10, 8.763382e-10, 8.753713e-10, 8.733474e-10, 8.737149e-10, 
    8.752016e-10, 8.785715e-10, 8.77428e-10, 8.803105e-10, 8.802454e-10, 
    8.834532e-10, 8.82007e-10, 8.873973e-10, 8.858657e-10, 8.902912e-10, 
    8.891784e-10, 8.902389e-10, 8.899174e-10, 8.90243e-10, 8.88611e-10, 
    8.893102e-10, 8.878741e-10, 8.822778e-10, 8.839227e-10, 8.790157e-10, 
    8.760634e-10, 8.741029e-10, 8.727111e-10, 8.729079e-10, 8.732829e-10, 
    8.752103e-10, 8.770223e-10, 8.78403e-10, 8.793263e-10, 8.802361e-10, 
    8.829882e-10, 8.844455e-10, 8.877067e-10, 8.871187e-10, 8.881152e-10, 
    8.890677e-10, 8.906661e-10, 8.904031e-10, 8.911071e-10, 8.880892e-10, 
    8.900949e-10, 8.867835e-10, 8.876893e-10, 8.804821e-10, 8.777366e-10, 
    8.765683e-10, 8.755465e-10, 8.730592e-10, 8.747768e-10, 8.740997e-10, 
    8.757108e-10, 8.767342e-10, 8.762281e-10, 8.793515e-10, 8.781373e-10, 
    8.845318e-10, 8.81778e-10, 8.889566e-10, 8.872394e-10, 8.893681e-10, 
    8.882821e-10, 8.901429e-10, 8.884682e-10, 8.913693e-10, 8.920008e-10, 
    8.915692e-10, 8.932272e-10, 8.883753e-10, 8.902387e-10, 8.762139e-10, 
    8.762964e-10, 8.76681e-10, 8.749901e-10, 8.748867e-10, 8.733372e-10, 
    8.747161e-10, 8.753031e-10, 8.767936e-10, 8.776749e-10, 8.785127e-10, 
    8.803543e-10, 8.824106e-10, 8.852856e-10, 8.873507e-10, 8.887346e-10, 
    8.878861e-10, 8.886352e-10, 8.877978e-10, 8.874053e-10, 8.917641e-10, 
    8.893167e-10, 8.929887e-10, 8.927857e-10, 8.911239e-10, 8.928085e-10, 
    8.763544e-10, 8.758794e-10, 8.742297e-10, 8.755207e-10, 8.731685e-10, 
    8.744851e-10, 8.75242e-10, 8.781624e-10, 8.788043e-10, 8.793989e-10, 
    8.805737e-10, 8.82081e-10, 8.847246e-10, 8.870241e-10, 8.891231e-10, 
    8.889693e-10, 8.890235e-10, 8.894922e-10, 8.88331e-10, 8.896828e-10, 
    8.899096e-10, 8.893166e-10, 8.927584e-10, 8.917753e-10, 8.927813e-10, 
    8.921412e-10, 8.760338e-10, 8.768331e-10, 8.764012e-10, 8.772132e-10, 
    8.766411e-10, 8.791848e-10, 8.799474e-10, 8.835149e-10, 8.820513e-10, 
    8.84381e-10, 8.822881e-10, 8.826589e-10, 8.844565e-10, 8.824013e-10, 
    8.868971e-10, 8.838489e-10, 8.895104e-10, 8.864668e-10, 8.897011e-10, 
    8.891141e-10, 8.900861e-10, 8.909565e-10, 8.920516e-10, 8.940714e-10, 
    8.936038e-10, 8.95293e-10, 8.780247e-10, 8.790609e-10, 8.7897e-10, 
    8.800545e-10, 8.808566e-10, 8.825949e-10, 8.85382e-10, 8.843341e-10, 
    8.86258e-10, 8.866441e-10, 8.837213e-10, 8.855158e-10, 8.797547e-10, 
    8.806855e-10, 8.801314e-10, 8.781063e-10, 8.845752e-10, 8.812558e-10, 
    8.873847e-10, 8.855872e-10, 8.908324e-10, 8.88224e-10, 8.933463e-10, 
    8.955346e-10, 8.975947e-10, 9.000004e-10, 8.796268e-10, 8.789227e-10, 
    8.801836e-10, 8.819275e-10, 8.83546e-10, 8.856968e-10, 8.85917e-10, 
    8.863198e-10, 8.873634e-10, 8.882406e-10, 8.86447e-10, 8.884605e-10, 
    8.809009e-10, 8.848634e-10, 8.786562e-10, 8.805254e-10, 8.818248e-10, 
    8.812551e-10, 8.842144e-10, 8.849116e-10, 8.877444e-10, 8.862803e-10, 
    8.949943e-10, 8.9114e-10, 9.018324e-10, 8.988455e-10, 8.786765e-10, 
    8.796245e-10, 8.829225e-10, 8.813535e-10, 8.858405e-10, 8.869445e-10, 
    8.878422e-10, 8.88989e-10, 8.891131e-10, 8.897925e-10, 8.88679e-10, 
    8.897486e-10, 8.857014e-10, 8.875103e-10, 8.825459e-10, 8.837543e-10, 
    8.831984e-10, 8.825886e-10, 8.844708e-10, 8.864751e-10, 8.865183e-10, 
    8.871608e-10, 8.889706e-10, 8.858588e-10, 8.954909e-10, 8.895429e-10, 
    8.80658e-10, 8.824829e-10, 8.827439e-10, 8.82037e-10, 8.868338e-10, 
    8.850961e-10, 8.89776e-10, 8.885115e-10, 8.905834e-10, 8.895539e-10, 
    8.894024e-10, 8.8808e-10, 8.872564e-10, 8.851757e-10, 8.834823e-10, 
    8.821396e-10, 8.824519e-10, 8.839268e-10, 8.865978e-10, 8.891241e-10, 
    8.885707e-10, 8.90426e-10, 8.855153e-10, 8.875745e-10, 8.867786e-10, 
    8.888539e-10, 8.843062e-10, 8.881778e-10, 8.833161e-10, 8.837426e-10, 
    8.850616e-10, 8.877139e-10, 8.883012e-10, 8.889275e-10, 8.885411e-10, 
    8.866657e-10, 8.863585e-10, 8.850296e-10, 8.846625e-10, 8.836498e-10, 
    8.828111e-10, 8.835773e-10, 8.843817e-10, 8.866666e-10, 8.88725e-10, 
    8.909687e-10, 8.91518e-10, 8.941378e-10, 8.920047e-10, 8.95524e-10, 
    8.925313e-10, 8.977117e-10, 8.884028e-10, 8.924439e-10, 8.851217e-10, 
    8.859109e-10, 8.873378e-10, 8.906104e-10, 8.888442e-10, 8.9091e-10, 
    8.863465e-10, 8.839776e-10, 8.833649e-10, 8.822212e-10, 8.833911e-10, 
    8.832959e-10, 8.844153e-10, 8.840557e-10, 8.867425e-10, 8.852993e-10, 
    8.893985e-10, 8.908938e-10, 8.951158e-10, 8.977029e-10, 9.003361e-10, 
    9.014983e-10, 9.01852e-10, 9.019999e-10 ;

 SOIL2C =
  5.784273, 5.784277, 5.784276, 5.78428, 5.784278, 5.784281, 5.784274, 
    5.784277, 5.784275, 5.784273, 5.784287, 5.78428, 5.784295, 5.78429, 
    5.784301, 5.784294, 5.784303, 5.784301, 5.784307, 5.784305, 5.784312, 
    5.784307, 5.784315, 5.78431, 5.784311, 5.784307, 5.784282, 5.784286, 
    5.784282, 5.784282, 5.784282, 5.784278, 5.784276, 5.784273, 5.784273, 
    5.784276, 5.784283, 5.78428, 5.784286, 5.784286, 5.784292, 5.784289, 
    5.784299, 5.784297, 5.784305, 5.784303, 5.784305, 5.784304, 5.784305, 
    5.784302, 5.784303, 5.7843, 5.78429, 5.784293, 5.784284, 5.784278, 
    5.784274, 5.784271, 5.784272, 5.784272, 5.784276, 5.78428, 5.784282, 
    5.784284, 5.784286, 5.784291, 5.784294, 5.7843, 5.784299, 5.784301, 
    5.784303, 5.784306, 5.784305, 5.784307, 5.784301, 5.784305, 5.784298, 
    5.7843, 5.784286, 5.784281, 5.784279, 5.784277, 5.784272, 5.784275, 
    5.784274, 5.784277, 5.784279, 5.784278, 5.784284, 5.784282, 5.784294, 
    5.784289, 5.784302, 5.784299, 5.784303, 5.784301, 5.784305, 5.784302, 
    5.784307, 5.784308, 5.784307, 5.784311, 5.784301, 5.784305, 5.784278, 
    5.784278, 5.784279, 5.784276, 5.784276, 5.784273, 5.784275, 5.784276, 
    5.784279, 5.784281, 5.784283, 5.784286, 5.78429, 5.784296, 5.784299, 
    5.784302, 5.7843, 5.784302, 5.7843, 5.784299, 5.784308, 5.784303, 
    5.78431, 5.78431, 5.784307, 5.78431, 5.784278, 5.784277, 5.784274, 
    5.784276, 5.784272, 5.784275, 5.784276, 5.784282, 5.784283, 5.784284, 
    5.784286, 5.784289, 5.784294, 5.784299, 5.784303, 5.784303, 5.784303, 
    5.784304, 5.784301, 5.784304, 5.784304, 5.784303, 5.78431, 5.784308, 
    5.78431, 5.784308, 5.784278, 5.784279, 5.784278, 5.78428, 5.784279, 
    5.784284, 5.784285, 5.784292, 5.784289, 5.784294, 5.78429, 5.78429, 
    5.784294, 5.78429, 5.784298, 5.784293, 5.784304, 5.784297, 5.784304, 
    5.784303, 5.784305, 5.784306, 5.784308, 5.784312, 5.784311, 5.784315, 
    5.784282, 5.784284, 5.784283, 5.784286, 5.784287, 5.78429, 5.784296, 
    5.784294, 5.784297, 5.784298, 5.784292, 5.784296, 5.784285, 5.784286, 
    5.784286, 5.784282, 5.784294, 5.784288, 5.784299, 5.784296, 5.784306, 
    5.784301, 5.784311, 5.784315, 5.784319, 5.784324, 5.784285, 5.784283, 
    5.784286, 5.784289, 5.784292, 5.784296, 5.784297, 5.784297, 5.784299, 
    5.784301, 5.784297, 5.784301, 5.784287, 5.784295, 5.784283, 5.784286, 
    5.784289, 5.784288, 5.784293, 5.784295, 5.7843, 5.784297, 5.784314, 
    5.784307, 5.784327, 5.784321, 5.784283, 5.784285, 5.784291, 5.784288, 
    5.784297, 5.784298, 5.7843, 5.784303, 5.784303, 5.784304, 5.784302, 
    5.784304, 5.784296, 5.7843, 5.78429, 5.784293, 5.784291, 5.78429, 
    5.784294, 5.784297, 5.784298, 5.784299, 5.784303, 5.784297, 5.784315, 
    5.784304, 5.784286, 5.78429, 5.784291, 5.784289, 5.784298, 5.784295, 
    5.784304, 5.784302, 5.784306, 5.784304, 5.784303, 5.784301, 5.784299, 
    5.784295, 5.784292, 5.784289, 5.78429, 5.784293, 5.784298, 5.784303, 
    5.784302, 5.784305, 5.784296, 5.7843, 5.784298, 5.784302, 5.784294, 
    5.784301, 5.784292, 5.784293, 5.784295, 5.7843, 5.784301, 5.784302, 
    5.784302, 5.784298, 5.784297, 5.784295, 5.784294, 5.784292, 5.784291, 
    5.784292, 5.784294, 5.784298, 5.784302, 5.784307, 5.784307, 5.784312, 
    5.784308, 5.784315, 5.784309, 5.784319, 5.784301, 5.784309, 5.784295, 
    5.784297, 5.784299, 5.784306, 5.784302, 5.784306, 5.784297, 5.784293, 
    5.784292, 5.784289, 5.784292, 5.784292, 5.784294, 5.784293, 5.784298, 
    5.784296, 5.784303, 5.784306, 5.784314, 5.784319, 5.784324, 5.784327, 
    5.784327, 5.784328 ;

 SOIL2C_TO_SOIL1C =
  1.302747e-09, 1.306316e-09, 1.305623e-09, 1.3085e-09, 1.306904e-09, 
    1.308788e-09, 1.303471e-09, 1.306458e-09, 1.304551e-09, 1.303069e-09, 
    1.314083e-09, 1.308629e-09, 1.319748e-09, 1.316271e-09, 1.325004e-09, 
    1.319207e-09, 1.326173e-09, 1.324838e-09, 1.328858e-09, 1.327706e-09, 
    1.332846e-09, 1.329389e-09, 1.335511e-09, 1.332021e-09, 1.332567e-09, 
    1.329275e-09, 1.309727e-09, 1.313404e-09, 1.309509e-09, 1.310034e-09, 
    1.309798e-09, 1.306937e-09, 1.305495e-09, 1.302475e-09, 1.303023e-09, 
    1.305241e-09, 1.310269e-09, 1.308563e-09, 1.312864e-09, 1.312767e-09, 
    1.317553e-09, 1.315395e-09, 1.323437e-09, 1.321152e-09, 1.327754e-09, 
    1.326094e-09, 1.327676e-09, 1.327197e-09, 1.327683e-09, 1.325248e-09, 
    1.326291e-09, 1.324148e-09, 1.315799e-09, 1.318253e-09, 1.310932e-09, 
    1.306527e-09, 1.303602e-09, 1.301526e-09, 1.301819e-09, 1.302379e-09, 
    1.305254e-09, 1.307958e-09, 1.310018e-09, 1.311395e-09, 1.312753e-09, 
    1.316859e-09, 1.319033e-09, 1.323899e-09, 1.323021e-09, 1.324508e-09, 
    1.325929e-09, 1.328314e-09, 1.327921e-09, 1.328972e-09, 1.324469e-09, 
    1.327461e-09, 1.322521e-09, 1.323873e-09, 1.31312e-09, 1.309024e-09, 
    1.30728e-09, 1.305756e-09, 1.302045e-09, 1.304608e-09, 1.303597e-09, 
    1.306001e-09, 1.307528e-09, 1.306773e-09, 1.311433e-09, 1.309621e-09, 
    1.319162e-09, 1.315053e-09, 1.325763e-09, 1.323201e-09, 1.326377e-09, 
    1.324757e-09, 1.327533e-09, 1.325035e-09, 1.329363e-09, 1.330305e-09, 
    1.329661e-09, 1.332135e-09, 1.324896e-09, 1.327676e-09, 1.306752e-09, 
    1.306875e-09, 1.307449e-09, 1.304926e-09, 1.304772e-09, 1.30246e-09, 
    1.304517e-09, 1.305393e-09, 1.307617e-09, 1.308932e-09, 1.310182e-09, 
    1.312929e-09, 1.315997e-09, 1.320286e-09, 1.323367e-09, 1.325432e-09, 
    1.324166e-09, 1.325284e-09, 1.324034e-09, 1.323449e-09, 1.329952e-09, 
    1.326301e-09, 1.331779e-09, 1.331476e-09, 1.328997e-09, 1.33151e-09, 
    1.306961e-09, 1.306253e-09, 1.303791e-09, 1.305718e-09, 1.302208e-09, 
    1.304172e-09, 1.305302e-09, 1.309659e-09, 1.310617e-09, 1.311504e-09, 
    1.313257e-09, 1.315505e-09, 1.319449e-09, 1.32288e-09, 1.326012e-09, 
    1.325782e-09, 1.325863e-09, 1.326562e-09, 1.32483e-09, 1.326847e-09, 
    1.327185e-09, 1.3263e-09, 1.331435e-09, 1.329968e-09, 1.331469e-09, 
    1.330514e-09, 1.306483e-09, 1.307676e-09, 1.307031e-09, 1.308243e-09, 
    1.307389e-09, 1.311184e-09, 1.312322e-09, 1.317645e-09, 1.315461e-09, 
    1.318937e-09, 1.315814e-09, 1.316367e-09, 1.319049e-09, 1.315983e-09, 
    1.322691e-09, 1.318143e-09, 1.32659e-09, 1.322049e-09, 1.326874e-09, 
    1.325998e-09, 1.327448e-09, 1.328747e-09, 1.330381e-09, 1.333394e-09, 
    1.332696e-09, 1.335216e-09, 1.309453e-09, 1.311e-09, 1.310864e-09, 
    1.312482e-09, 1.313678e-09, 1.316272e-09, 1.32043e-09, 1.318867e-09, 
    1.321737e-09, 1.322313e-09, 1.317953e-09, 1.32063e-09, 1.312034e-09, 
    1.313423e-09, 1.312597e-09, 1.309575e-09, 1.319227e-09, 1.314274e-09, 
    1.323418e-09, 1.320736e-09, 1.328562e-09, 1.32467e-09, 1.332312e-09, 
    1.335577e-09, 1.33865e-09, 1.342239e-09, 1.311844e-09, 1.310793e-09, 
    1.312675e-09, 1.315276e-09, 1.317691e-09, 1.3209e-09, 1.321228e-09, 
    1.321829e-09, 1.323386e-09, 1.324695e-09, 1.322019e-09, 1.325023e-09, 
    1.313745e-09, 1.319656e-09, 1.310396e-09, 1.313184e-09, 1.315123e-09, 
    1.314273e-09, 1.318688e-09, 1.319729e-09, 1.323955e-09, 1.32177e-09, 
    1.334771e-09, 1.329021e-09, 1.344972e-09, 1.340516e-09, 1.310426e-09, 
    1.31184e-09, 1.316761e-09, 1.31442e-09, 1.321114e-09, 1.322761e-09, 
    1.324101e-09, 1.325812e-09, 1.325997e-09, 1.32701e-09, 1.325349e-09, 
    1.326945e-09, 1.320907e-09, 1.323605e-09, 1.316199e-09, 1.318002e-09, 
    1.317172e-09, 1.316263e-09, 1.319071e-09, 1.322061e-09, 1.322126e-09, 
    1.323084e-09, 1.325784e-09, 1.321142e-09, 1.335512e-09, 1.326638e-09, 
    1.313382e-09, 1.316105e-09, 1.316494e-09, 1.31544e-09, 1.322596e-09, 
    1.320004e-09, 1.326986e-09, 1.325099e-09, 1.32819e-09, 1.326654e-09, 
    1.326428e-09, 1.324455e-09, 1.323227e-09, 1.320122e-09, 1.317596e-09, 
    1.315593e-09, 1.316059e-09, 1.318259e-09, 1.322244e-09, 1.326013e-09, 
    1.325188e-09, 1.327955e-09, 1.320629e-09, 1.323701e-09, 1.322514e-09, 
    1.32561e-09, 1.318825e-09, 1.324601e-09, 1.317348e-09, 1.317984e-09, 
    1.319952e-09, 1.323909e-09, 1.324786e-09, 1.32572e-09, 1.325143e-09, 
    1.322345e-09, 1.321887e-09, 1.319904e-09, 1.319357e-09, 1.317846e-09, 
    1.316595e-09, 1.317738e-09, 1.318938e-09, 1.322347e-09, 1.325418e-09, 
    1.328765e-09, 1.329585e-09, 1.333493e-09, 1.330311e-09, 1.335561e-09, 
    1.331096e-09, 1.338825e-09, 1.324937e-09, 1.330966e-09, 1.320042e-09, 
    1.321219e-09, 1.323348e-09, 1.328231e-09, 1.325596e-09, 1.328678e-09, 
    1.321869e-09, 1.318335e-09, 1.317421e-09, 1.315714e-09, 1.31746e-09, 
    1.317318e-09, 1.318988e-09, 1.318451e-09, 1.32246e-09, 1.320307e-09, 
    1.326423e-09, 1.328653e-09, 1.334952e-09, 1.338812e-09, 1.34274e-09, 
    1.344474e-09, 1.345002e-09, 1.345222e-09 ;

 SOIL2C_TO_SOIL3C =
  9.305338e-11, 9.330831e-11, 9.325876e-11, 9.346431e-11, 9.335031e-11, 
    9.348489e-11, 9.310509e-11, 9.33184e-11, 9.318225e-11, 9.307636e-11, 
    9.386304e-11, 9.347349e-11, 9.42677e-11, 9.401935e-11, 9.464315e-11, 
    9.422904e-11, 9.472664e-11, 9.463125e-11, 9.491842e-11, 9.483616e-11, 
    9.520329e-11, 9.495639e-11, 9.539361e-11, 9.514436e-11, 9.518333e-11, 
    9.494824e-11, 9.355194e-11, 9.381454e-11, 9.353637e-11, 9.357382e-11, 
    9.355702e-11, 9.335265e-11, 9.324962e-11, 9.303392e-11, 9.307309e-11, 
    9.323153e-11, 9.359066e-11, 9.34688e-11, 9.377598e-11, 9.376905e-11, 
    9.41109e-11, 9.395678e-11, 9.453121e-11, 9.436799e-11, 9.483959e-11, 
    9.472101e-11, 9.483402e-11, 9.479976e-11, 9.483447e-11, 9.466054e-11, 
    9.473506e-11, 9.458202e-11, 9.398564e-11, 9.416093e-11, 9.3638e-11, 
    9.332338e-11, 9.311443e-11, 9.296611e-11, 9.298708e-11, 9.302705e-11, 
    9.323246e-11, 9.342557e-11, 9.35727e-11, 9.36711e-11, 9.376806e-11, 
    9.406135e-11, 9.421664e-11, 9.456418e-11, 9.450151e-11, 9.460771e-11, 
    9.470921e-11, 9.487955e-11, 9.485152e-11, 9.492655e-11, 9.460494e-11, 
    9.481868e-11, 9.44658e-11, 9.456232e-11, 9.379427e-11, 9.350168e-11, 
    9.337717e-11, 9.326828e-11, 9.300321e-11, 9.318626e-11, 9.31141e-11, 
    9.328579e-11, 9.339486e-11, 9.334093e-11, 9.367379e-11, 9.354439e-11, 
    9.422584e-11, 9.393238e-11, 9.469737e-11, 9.451438e-11, 9.474124e-11, 
    9.462549e-11, 9.482379e-11, 9.464533e-11, 9.495448e-11, 9.502178e-11, 
    9.497579e-11, 9.515247e-11, 9.463543e-11, 9.483401e-11, 9.333941e-11, 
    9.33482e-11, 9.338919e-11, 9.320899e-11, 9.319797e-11, 9.303284e-11, 
    9.317979e-11, 9.324234e-11, 9.340119e-11, 9.349511e-11, 9.358439e-11, 
    9.378066e-11, 9.399979e-11, 9.430617e-11, 9.452624e-11, 9.467372e-11, 
    9.45833e-11, 9.466313e-11, 9.457388e-11, 9.453206e-11, 9.499655e-11, 
    9.473575e-11, 9.512706e-11, 9.510542e-11, 9.492833e-11, 9.510785e-11, 
    9.335438e-11, 9.330376e-11, 9.312795e-11, 9.326554e-11, 9.301486e-11, 
    9.315516e-11, 9.323583e-11, 9.354706e-11, 9.361547e-11, 9.367884e-11, 
    9.380404e-11, 9.396467e-11, 9.424638e-11, 9.449144e-11, 9.471512e-11, 
    9.469873e-11, 9.470451e-11, 9.475445e-11, 9.463071e-11, 9.477476e-11, 
    9.479893e-11, 9.473573e-11, 9.510252e-11, 9.499775e-11, 9.510495e-11, 
    9.503675e-11, 9.332022e-11, 9.340539e-11, 9.335937e-11, 9.344591e-11, 
    9.338493e-11, 9.365602e-11, 9.373729e-11, 9.411748e-11, 9.39615e-11, 
    9.420977e-11, 9.398674e-11, 9.402625e-11, 9.421781e-11, 9.399879e-11, 
    9.44779e-11, 9.415307e-11, 9.475639e-11, 9.443205e-11, 9.477671e-11, 
    9.471415e-11, 9.481774e-11, 9.491049e-11, 9.502719e-11, 9.524243e-11, 
    9.51926e-11, 9.53726e-11, 9.353238e-11, 9.364282e-11, 9.363312e-11, 
    9.374871e-11, 9.383418e-11, 9.401942e-11, 9.431644e-11, 9.420478e-11, 
    9.44098e-11, 9.445095e-11, 9.413947e-11, 9.43307e-11, 9.371675e-11, 
    9.381594e-11, 9.375691e-11, 9.354108e-11, 9.423047e-11, 9.387672e-11, 
    9.452987e-11, 9.433831e-11, 9.489726e-11, 9.461931e-11, 9.516516e-11, 
    9.539835e-11, 9.561788e-11, 9.587423e-11, 9.370312e-11, 9.362808e-11, 
    9.376246e-11, 9.394831e-11, 9.412079e-11, 9.434999e-11, 9.437346e-11, 
    9.441638e-11, 9.452759e-11, 9.462107e-11, 9.442993e-11, 9.464451e-11, 
    9.38389e-11, 9.426118e-11, 9.359969e-11, 9.379889e-11, 9.393736e-11, 
    9.387665e-11, 9.419202e-11, 9.426632e-11, 9.456819e-11, 9.441217e-11, 
    9.534078e-11, 9.493005e-11, 9.606946e-11, 9.575116e-11, 9.360186e-11, 
    9.370287e-11, 9.405434e-11, 9.388713e-11, 9.436531e-11, 9.448296e-11, 
    9.457862e-11, 9.470084e-11, 9.471405e-11, 9.478646e-11, 9.466779e-11, 
    9.478178e-11, 9.435049e-11, 9.454325e-11, 9.401421e-11, 9.414299e-11, 
    9.408375e-11, 9.401876e-11, 9.421933e-11, 9.443293e-11, 9.443754e-11, 
    9.450601e-11, 9.469886e-11, 9.436725e-11, 9.539369e-11, 9.475985e-11, 
    9.381302e-11, 9.400749e-11, 9.403531e-11, 9.395998e-11, 9.447116e-11, 
    9.428597e-11, 9.47847e-11, 9.464995e-11, 9.487074e-11, 9.476103e-11, 
    9.474488e-11, 9.460396e-11, 9.45162e-11, 9.429445e-11, 9.4114e-11, 
    9.397091e-11, 9.400419e-11, 9.416137e-11, 9.444601e-11, 9.471522e-11, 
    9.465626e-11, 9.485396e-11, 9.433065e-11, 9.45501e-11, 9.446528e-11, 
    9.468644e-11, 9.420181e-11, 9.461439e-11, 9.409629e-11, 9.414174e-11, 
    9.42823e-11, 9.456495e-11, 9.462753e-11, 9.469427e-11, 9.46531e-11, 
    9.445324e-11, 9.442051e-11, 9.427889e-11, 9.423976e-11, 9.413185e-11, 
    9.404247e-11, 9.412412e-11, 9.420986e-11, 9.445334e-11, 9.46727e-11, 
    9.49118e-11, 9.497033e-11, 9.52495e-11, 9.50222e-11, 9.539722e-11, 
    9.507831e-11, 9.563034e-11, 9.463836e-11, 9.5069e-11, 9.428871e-11, 
    9.437281e-11, 9.452487e-11, 9.487362e-11, 9.46854e-11, 9.490553e-11, 
    9.441923e-11, 9.416678e-11, 9.410149e-11, 9.397961e-11, 9.410428e-11, 
    9.409414e-11, 9.421343e-11, 9.41751e-11, 9.446142e-11, 9.430764e-11, 
    9.474446e-11, 9.490381e-11, 9.535372e-11, 9.56294e-11, 9.591001e-11, 
    9.603385e-11, 9.607154e-11, 9.60873e-11 ;

 SOIL2C_vr =
  20.00613, 20.00614, 20.00614, 20.00615, 20.00614, 20.00615, 20.00613, 
    20.00614, 20.00613, 20.00613, 20.00618, 20.00615, 20.0062, 20.00619, 
    20.00622, 20.0062, 20.00623, 20.00622, 20.00624, 20.00624, 20.00626, 
    20.00624, 20.00627, 20.00625, 20.00626, 20.00624, 20.00616, 20.00617, 
    20.00616, 20.00616, 20.00616, 20.00614, 20.00614, 20.00612, 20.00613, 
    20.00614, 20.00616, 20.00615, 20.00617, 20.00617, 20.00619, 20.00618, 
    20.00622, 20.00621, 20.00624, 20.00623, 20.00624, 20.00623, 20.00624, 
    20.00622, 20.00623, 20.00622, 20.00618, 20.00619, 20.00616, 20.00614, 
    20.00613, 20.00612, 20.00612, 20.00612, 20.00614, 20.00615, 20.00616, 
    20.00616, 20.00617, 20.00619, 20.0062, 20.00622, 20.00621, 20.00622, 
    20.00623, 20.00624, 20.00624, 20.00624, 20.00622, 20.00624, 20.00621, 
    20.00622, 20.00617, 20.00615, 20.00615, 20.00614, 20.00612, 20.00613, 
    20.00613, 20.00614, 20.00615, 20.00614, 20.00616, 20.00616, 20.0062, 
    20.00618, 20.00623, 20.00622, 20.00623, 20.00622, 20.00624, 20.00622, 
    20.00624, 20.00625, 20.00624, 20.00625, 20.00622, 20.00624, 20.00614, 
    20.00614, 20.00615, 20.00614, 20.00613, 20.00612, 20.00613, 20.00614, 
    20.00615, 20.00615, 20.00616, 20.00617, 20.00618, 20.0062, 20.00622, 
    20.00623, 20.00622, 20.00623, 20.00622, 20.00622, 20.00624, 20.00623, 
    20.00625, 20.00625, 20.00624, 20.00625, 20.00614, 20.00614, 20.00613, 
    20.00614, 20.00612, 20.00613, 20.00614, 20.00616, 20.00616, 20.00616, 
    20.00617, 20.00618, 20.0062, 20.00621, 20.00623, 20.00623, 20.00623, 
    20.00623, 20.00622, 20.00623, 20.00623, 20.00623, 20.00625, 20.00624, 
    20.00625, 20.00625, 20.00614, 20.00615, 20.00614, 20.00615, 20.00615, 
    20.00616, 20.00617, 20.00619, 20.00618, 20.0062, 20.00618, 20.00619, 
    20.0062, 20.00618, 20.00621, 20.00619, 20.00623, 20.00621, 20.00623, 
    20.00623, 20.00624, 20.00624, 20.00625, 20.00626, 20.00626, 20.00627, 
    20.00616, 20.00616, 20.00616, 20.00617, 20.00617, 20.00619, 20.0062, 
    20.0062, 20.00621, 20.00621, 20.00619, 20.0062, 20.00617, 20.00617, 
    20.00617, 20.00616, 20.0062, 20.00618, 20.00622, 20.0062, 20.00624, 
    20.00622, 20.00626, 20.00627, 20.00628, 20.0063, 20.00617, 20.00616, 
    20.00617, 20.00618, 20.00619, 20.0062, 20.00621, 20.00621, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00617, 20.0062, 20.00616, 20.00617, 
    20.00618, 20.00618, 20.0062, 20.0062, 20.00622, 20.00621, 20.00627, 
    20.00624, 20.00631, 20.00629, 20.00616, 20.00617, 20.00619, 20.00618, 
    20.00621, 20.00621, 20.00622, 20.00623, 20.00623, 20.00623, 20.00623, 
    20.00623, 20.0062, 20.00622, 20.00619, 20.00619, 20.00619, 20.00619, 
    20.0062, 20.00621, 20.00621, 20.00621, 20.00623, 20.00621, 20.00627, 
    20.00623, 20.00617, 20.00618, 20.00619, 20.00618, 20.00621, 20.0062, 
    20.00623, 20.00622, 20.00624, 20.00623, 20.00623, 20.00622, 20.00622, 
    20.0062, 20.00619, 20.00618, 20.00618, 20.00619, 20.00621, 20.00623, 
    20.00622, 20.00624, 20.0062, 20.00622, 20.00621, 20.00623, 20.0062, 
    20.00622, 20.00619, 20.00619, 20.0062, 20.00622, 20.00622, 20.00623, 
    20.00622, 20.00621, 20.00621, 20.0062, 20.0062, 20.00619, 20.00619, 
    20.00619, 20.0062, 20.00621, 20.00623, 20.00624, 20.00624, 20.00626, 
    20.00625, 20.00627, 20.00625, 20.00628, 20.00622, 20.00625, 20.0062, 
    20.00621, 20.00622, 20.00624, 20.00623, 20.00624, 20.00621, 20.0062, 
    20.00619, 20.00618, 20.00619, 20.00619, 20.0062, 20.0062, 20.00621, 
    20.0062, 20.00623, 20.00624, 20.00627, 20.00628, 20.0063, 20.00631, 
    20.00631, 20.00631,
  20.00632, 20.00634, 20.00633, 20.00635, 20.00634, 20.00635, 20.00632, 
    20.00634, 20.00633, 20.00632, 20.00637, 20.00635, 20.0064, 20.00638, 
    20.00642, 20.0064, 20.00643, 20.00642, 20.00644, 20.00644, 20.00646, 
    20.00644, 20.00647, 20.00646, 20.00646, 20.00644, 20.00635, 20.00637, 
    20.00635, 20.00635, 20.00635, 20.00634, 20.00633, 20.00632, 20.00632, 
    20.00633, 20.00636, 20.00635, 20.00637, 20.00637, 20.00639, 20.00638, 
    20.00642, 20.0064, 20.00644, 20.00643, 20.00644, 20.00643, 20.00644, 
    20.00642, 20.00643, 20.00642, 20.00638, 20.00639, 20.00636, 20.00634, 
    20.00632, 20.00631, 20.00632, 20.00632, 20.00633, 20.00634, 20.00635, 
    20.00636, 20.00637, 20.00639, 20.0064, 20.00642, 20.00641, 20.00642, 
    20.00643, 20.00644, 20.00644, 20.00644, 20.00642, 20.00644, 20.00641, 
    20.00642, 20.00637, 20.00635, 20.00634, 20.00633, 20.00632, 20.00633, 
    20.00632, 20.00633, 20.00634, 20.00634, 20.00636, 20.00635, 20.0064, 
    20.00638, 20.00643, 20.00641, 20.00643, 20.00642, 20.00644, 20.00642, 
    20.00644, 20.00645, 20.00644, 20.00646, 20.00642, 20.00644, 20.00634, 
    20.00634, 20.00634, 20.00633, 20.00633, 20.00632, 20.00633, 20.00633, 
    20.00634, 20.00635, 20.00635, 20.00637, 20.00638, 20.0064, 20.00642, 
    20.00643, 20.00642, 20.00642, 20.00642, 20.00642, 20.00645, 20.00643, 
    20.00645, 20.00645, 20.00644, 20.00645, 20.00634, 20.00634, 20.00632, 
    20.00633, 20.00632, 20.00633, 20.00633, 20.00635, 20.00636, 20.00636, 
    20.00637, 20.00638, 20.0064, 20.00641, 20.00643, 20.00643, 20.00643, 
    20.00643, 20.00642, 20.00643, 20.00643, 20.00643, 20.00645, 20.00645, 
    20.00645, 20.00645, 20.00634, 20.00634, 20.00634, 20.00635, 20.00634, 
    20.00636, 20.00636, 20.00639, 20.00638, 20.0064, 20.00638, 20.00638, 
    20.0064, 20.00638, 20.00641, 20.00639, 20.00643, 20.00641, 20.00643, 
    20.00643, 20.00644, 20.00644, 20.00645, 20.00646, 20.00646, 20.00647, 
    20.00635, 20.00636, 20.00636, 20.00636, 20.00637, 20.00638, 20.0064, 
    20.0064, 20.00641, 20.00641, 20.00639, 20.0064, 20.00636, 20.00637, 
    20.00636, 20.00635, 20.0064, 20.00637, 20.00642, 20.0064, 20.00644, 
    20.00642, 20.00646, 20.00647, 20.00649, 20.0065, 20.00636, 20.00636, 
    20.00637, 20.00638, 20.00639, 20.0064, 20.0064, 20.00641, 20.00642, 
    20.00642, 20.00641, 20.00642, 20.00637, 20.0064, 20.00636, 20.00637, 
    20.00638, 20.00637, 20.00639, 20.0064, 20.00642, 20.00641, 20.00647, 
    20.00644, 20.00652, 20.00649, 20.00636, 20.00636, 20.00639, 20.00637, 
    20.0064, 20.00641, 20.00642, 20.00643, 20.00643, 20.00643, 20.00643, 
    20.00643, 20.0064, 20.00642, 20.00638, 20.00639, 20.00639, 20.00638, 
    20.0064, 20.00641, 20.00641, 20.00641, 20.00643, 20.0064, 20.00647, 
    20.00643, 20.00637, 20.00638, 20.00638, 20.00638, 20.00641, 20.0064, 
    20.00643, 20.00642, 20.00644, 20.00643, 20.00643, 20.00642, 20.00641, 
    20.0064, 20.00639, 20.00638, 20.00638, 20.00639, 20.00641, 20.00643, 
    20.00642, 20.00644, 20.0064, 20.00642, 20.00641, 20.00643, 20.0064, 
    20.00642, 20.00639, 20.00639, 20.0064, 20.00642, 20.00642, 20.00643, 
    20.00642, 20.00641, 20.00641, 20.0064, 20.0064, 20.00639, 20.00638, 
    20.00639, 20.0064, 20.00641, 20.00643, 20.00644, 20.00644, 20.00646, 
    20.00645, 20.00647, 20.00645, 20.00649, 20.00642, 20.00645, 20.0064, 
    20.0064, 20.00642, 20.00644, 20.00643, 20.00644, 20.00641, 20.00639, 
    20.00639, 20.00638, 20.00639, 20.00639, 20.0064, 20.00639, 20.00641, 
    20.0064, 20.00643, 20.00644, 20.00647, 20.00649, 20.00651, 20.00651, 
    20.00652, 20.00652,
  20.00634, 20.00636, 20.00635, 20.00637, 20.00636, 20.00637, 20.00634, 
    20.00636, 20.00635, 20.00634, 20.00639, 20.00637, 20.00642, 20.0064, 
    20.00644, 20.00642, 20.00645, 20.00644, 20.00646, 20.00646, 20.00648, 
    20.00647, 20.00649, 20.00648, 20.00648, 20.00647, 20.00637, 20.00639, 
    20.00637, 20.00637, 20.00637, 20.00636, 20.00635, 20.00634, 20.00634, 
    20.00635, 20.00638, 20.00637, 20.00639, 20.00639, 20.00641, 20.0064, 
    20.00644, 20.00643, 20.00646, 20.00645, 20.00646, 20.00646, 20.00646, 
    20.00645, 20.00645, 20.00644, 20.0064, 20.00641, 20.00638, 20.00636, 
    20.00634, 20.00633, 20.00634, 20.00634, 20.00635, 20.00636, 20.00637, 
    20.00638, 20.00639, 20.00641, 20.00642, 20.00644, 20.00644, 20.00644, 
    20.00645, 20.00646, 20.00646, 20.00646, 20.00644, 20.00646, 20.00643, 
    20.00644, 20.00639, 20.00637, 20.00636, 20.00636, 20.00634, 20.00635, 
    20.00634, 20.00636, 20.00636, 20.00636, 20.00638, 20.00637, 20.00642, 
    20.0064, 20.00645, 20.00644, 20.00645, 20.00644, 20.00646, 20.00644, 
    20.00647, 20.00647, 20.00647, 20.00648, 20.00644, 20.00646, 20.00636, 
    20.00636, 20.00636, 20.00635, 20.00635, 20.00634, 20.00635, 20.00635, 
    20.00636, 20.00637, 20.00638, 20.00639, 20.0064, 20.00642, 20.00644, 
    20.00645, 20.00644, 20.00645, 20.00644, 20.00644, 20.00647, 20.00645, 
    20.00648, 20.00648, 20.00646, 20.00648, 20.00636, 20.00636, 20.00635, 
    20.00636, 20.00634, 20.00635, 20.00635, 20.00637, 20.00638, 20.00638, 
    20.00639, 20.0064, 20.00642, 20.00644, 20.00645, 20.00645, 20.00645, 
    20.00645, 20.00644, 20.00645, 20.00646, 20.00645, 20.00648, 20.00647, 
    20.00648, 20.00647, 20.00636, 20.00636, 20.00636, 20.00637, 20.00636, 
    20.00638, 20.00639, 20.00641, 20.0064, 20.00642, 20.0064, 20.0064, 
    20.00642, 20.0064, 20.00644, 20.00641, 20.00645, 20.00643, 20.00645, 
    20.00645, 20.00646, 20.00646, 20.00647, 20.00648, 20.00648, 20.00649, 
    20.00637, 20.00638, 20.00638, 20.00639, 20.00639, 20.0064, 20.00642, 
    20.00642, 20.00643, 20.00643, 20.00641, 20.00642, 20.00638, 20.00639, 
    20.00639, 20.00637, 20.00642, 20.0064, 20.00644, 20.00643, 20.00646, 
    20.00644, 20.00648, 20.00649, 20.00651, 20.00653, 20.00638, 20.00638, 
    20.00639, 20.0064, 20.00641, 20.00643, 20.00643, 20.00643, 20.00644, 
    20.00644, 20.00643, 20.00644, 20.00639, 20.00642, 20.00638, 20.00639, 
    20.0064, 20.0064, 20.00642, 20.00642, 20.00644, 20.00643, 20.00649, 
    20.00646, 20.00654, 20.00652, 20.00638, 20.00638, 20.00641, 20.0064, 
    20.00643, 20.00644, 20.00644, 20.00645, 20.00645, 20.00645, 20.00645, 
    20.00645, 20.00643, 20.00644, 20.0064, 20.00641, 20.00641, 20.0064, 
    20.00642, 20.00643, 20.00643, 20.00644, 20.00645, 20.00643, 20.00649, 
    20.00645, 20.00639, 20.0064, 20.0064, 20.0064, 20.00643, 20.00642, 
    20.00645, 20.00645, 20.00646, 20.00645, 20.00645, 20.00644, 20.00644, 
    20.00642, 20.00641, 20.0064, 20.0064, 20.00641, 20.00643, 20.00645, 
    20.00645, 20.00646, 20.00642, 20.00644, 20.00643, 20.00645, 20.00642, 
    20.00644, 20.00641, 20.00641, 20.00642, 20.00644, 20.00644, 20.00645, 
    20.00645, 20.00643, 20.00643, 20.00642, 20.00642, 20.00641, 20.0064, 
    20.00641, 20.00642, 20.00643, 20.00645, 20.00646, 20.00647, 20.00648, 
    20.00647, 20.00649, 20.00647, 20.00651, 20.00644, 20.00647, 20.00642, 
    20.00643, 20.00644, 20.00646, 20.00645, 20.00646, 20.00643, 20.00641, 
    20.00641, 20.0064, 20.00641, 20.00641, 20.00642, 20.00641, 20.00643, 
    20.00642, 20.00645, 20.00646, 20.00649, 20.00651, 20.00653, 20.00654, 
    20.00654, 20.00654,
  20.00615, 20.00616, 20.00616, 20.00617, 20.00617, 20.00617, 20.00615, 
    20.00616, 20.00616, 20.00615, 20.0062, 20.00617, 20.00623, 20.00621, 
    20.00625, 20.00622, 20.00626, 20.00625, 20.00627, 20.00626, 20.00629, 
    20.00627, 20.0063, 20.00628, 20.00629, 20.00627, 20.00618, 20.0062, 
    20.00618, 20.00618, 20.00618, 20.00617, 20.00616, 20.00615, 20.00615, 
    20.00616, 20.00618, 20.00617, 20.00619, 20.00619, 20.00622, 20.00621, 
    20.00624, 20.00623, 20.00626, 20.00626, 20.00626, 20.00626, 20.00626, 
    20.00625, 20.00626, 20.00625, 20.00621, 20.00622, 20.00619, 20.00616, 
    20.00615, 20.00614, 20.00614, 20.00615, 20.00616, 20.00617, 20.00618, 
    20.00619, 20.00619, 20.00621, 20.00622, 20.00624, 20.00624, 20.00625, 
    20.00625, 20.00627, 20.00626, 20.00627, 20.00625, 20.00626, 20.00624, 
    20.00624, 20.0062, 20.00618, 20.00617, 20.00616, 20.00614, 20.00616, 
    20.00615, 20.00616, 20.00617, 20.00616, 20.00619, 20.00618, 20.00622, 
    20.0062, 20.00625, 20.00624, 20.00626, 20.00625, 20.00626, 20.00625, 
    20.00627, 20.00628, 20.00627, 20.00628, 20.00625, 20.00626, 20.00616, 
    20.00617, 20.00617, 20.00616, 20.00616, 20.00615, 20.00616, 20.00616, 
    20.00617, 20.00618, 20.00618, 20.0062, 20.00621, 20.00623, 20.00624, 
    20.00625, 20.00625, 20.00625, 20.00625, 20.00624, 20.00627, 20.00626, 
    20.00628, 20.00628, 20.00627, 20.00628, 20.00617, 20.00616, 20.00615, 
    20.00616, 20.00614, 20.00615, 20.00616, 20.00618, 20.00618, 20.00619, 
    20.0062, 20.00621, 20.00623, 20.00624, 20.00626, 20.00625, 20.00625, 
    20.00626, 20.00625, 20.00626, 20.00626, 20.00626, 20.00628, 20.00627, 
    20.00628, 20.00628, 20.00616, 20.00617, 20.00617, 20.00617, 20.00617, 
    20.00619, 20.00619, 20.00622, 20.00621, 20.00622, 20.00621, 20.00621, 
    20.00622, 20.00621, 20.00624, 20.00622, 20.00626, 20.00624, 20.00626, 
    20.00626, 20.00626, 20.00627, 20.00628, 20.00629, 20.00629, 20.0063, 
    20.00618, 20.00619, 20.00618, 20.00619, 20.0062, 20.00621, 20.00623, 
    20.00622, 20.00624, 20.00624, 20.00622, 20.00623, 20.00619, 20.0062, 
    20.00619, 20.00618, 20.00622, 20.0062, 20.00624, 20.00623, 20.00627, 
    20.00625, 20.00628, 20.0063, 20.00631, 20.00633, 20.00619, 20.00618, 
    20.00619, 20.0062, 20.00622, 20.00623, 20.00623, 20.00624, 20.00624, 
    20.00625, 20.00624, 20.00625, 20.0062, 20.00623, 20.00618, 20.0062, 
    20.0062, 20.0062, 20.00622, 20.00623, 20.00625, 20.00624, 20.0063, 
    20.00627, 20.00634, 20.00632, 20.00618, 20.00619, 20.00621, 20.0062, 
    20.00623, 20.00624, 20.00625, 20.00625, 20.00626, 20.00626, 20.00625, 
    20.00626, 20.00623, 20.00624, 20.00621, 20.00622, 20.00621, 20.00621, 
    20.00622, 20.00624, 20.00624, 20.00624, 20.00625, 20.00623, 20.0063, 
    20.00626, 20.0062, 20.00621, 20.00621, 20.00621, 20.00624, 20.00623, 
    20.00626, 20.00625, 20.00627, 20.00626, 20.00626, 20.00625, 20.00624, 
    20.00623, 20.00622, 20.00621, 20.00621, 20.00622, 20.00624, 20.00626, 
    20.00625, 20.00626, 20.00623, 20.00624, 20.00624, 20.00625, 20.00622, 
    20.00625, 20.00621, 20.00622, 20.00623, 20.00624, 20.00625, 20.00625, 
    20.00625, 20.00624, 20.00624, 20.00623, 20.00622, 20.00622, 20.00621, 
    20.00622, 20.00622, 20.00624, 20.00625, 20.00627, 20.00627, 20.00629, 
    20.00628, 20.0063, 20.00628, 20.00632, 20.00625, 20.00628, 20.00623, 
    20.00623, 20.00624, 20.00627, 20.00625, 20.00627, 20.00624, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00621, 20.00622, 20.00622, 20.00624, 
    20.00623, 20.00626, 20.00627, 20.0063, 20.00632, 20.00633, 20.00634, 
    20.00634, 20.00635,
  20.00526, 20.00528, 20.00527, 20.00529, 20.00528, 20.00529, 20.00526, 
    20.00528, 20.00527, 20.00526, 20.00531, 20.00529, 20.00533, 20.00532, 
    20.00535, 20.00533, 20.00536, 20.00535, 20.00537, 20.00537, 20.00539, 
    20.00537, 20.0054, 20.00538, 20.00538, 20.00537, 20.00529, 20.00531, 
    20.00529, 20.00529, 20.00529, 20.00528, 20.00527, 20.00526, 20.00526, 
    20.00527, 20.00529, 20.00529, 20.0053, 20.0053, 20.00532, 20.00531, 
    20.00535, 20.00534, 20.00537, 20.00536, 20.00537, 20.00536, 20.00537, 
    20.00536, 20.00536, 20.00535, 20.00532, 20.00533, 20.00529, 20.00528, 
    20.00526, 20.00526, 20.00526, 20.00526, 20.00527, 20.00528, 20.00529, 
    20.0053, 20.0053, 20.00532, 20.00533, 20.00535, 20.00535, 20.00535, 
    20.00536, 20.00537, 20.00537, 20.00537, 20.00535, 20.00536, 20.00534, 
    20.00535, 20.0053, 20.00529, 20.00528, 20.00527, 20.00526, 20.00527, 
    20.00526, 20.00528, 20.00528, 20.00528, 20.0053, 20.00529, 20.00533, 
    20.00531, 20.00536, 20.00535, 20.00536, 20.00535, 20.00537, 20.00535, 
    20.00537, 20.00538, 20.00537, 20.00538, 20.00535, 20.00537, 20.00528, 
    20.00528, 20.00528, 20.00527, 20.00527, 20.00526, 20.00527, 20.00527, 
    20.00528, 20.00529, 20.00529, 20.0053, 20.00532, 20.00533, 20.00535, 
    20.00536, 20.00535, 20.00536, 20.00535, 20.00535, 20.00537, 20.00536, 
    20.00538, 20.00538, 20.00537, 20.00538, 20.00528, 20.00528, 20.00527, 
    20.00527, 20.00526, 20.00527, 20.00527, 20.00529, 20.00529, 20.0053, 
    20.0053, 20.00531, 20.00533, 20.00534, 20.00536, 20.00536, 20.00536, 
    20.00536, 20.00535, 20.00536, 20.00536, 20.00536, 20.00538, 20.00537, 
    20.00538, 20.00538, 20.00528, 20.00528, 20.00528, 20.00528, 20.00528, 
    20.0053, 20.0053, 20.00532, 20.00531, 20.00533, 20.00532, 20.00532, 
    20.00533, 20.00532, 20.00534, 20.00533, 20.00536, 20.00534, 20.00536, 
    20.00536, 20.00536, 20.00537, 20.00538, 20.00539, 20.00539, 20.0054, 
    20.00529, 20.00529, 20.00529, 20.0053, 20.00531, 20.00532, 20.00533, 
    20.00533, 20.00534, 20.00534, 20.00533, 20.00533, 20.0053, 20.00531, 
    20.0053, 20.00529, 20.00533, 20.00531, 20.00535, 20.00534, 20.00537, 
    20.00535, 20.00538, 20.0054, 20.00541, 20.00543, 20.0053, 20.00529, 
    20.0053, 20.00531, 20.00532, 20.00534, 20.00534, 20.00534, 20.00535, 
    20.00535, 20.00534, 20.00535, 20.00531, 20.00533, 20.00529, 20.0053, 
    20.00531, 20.00531, 20.00533, 20.00533, 20.00535, 20.00534, 20.00539, 
    20.00537, 20.00544, 20.00542, 20.00529, 20.0053, 20.00532, 20.00531, 
    20.00534, 20.00534, 20.00535, 20.00536, 20.00536, 20.00536, 20.00536, 
    20.00536, 20.00534, 20.00535, 20.00532, 20.00533, 20.00532, 20.00532, 
    20.00533, 20.00534, 20.00534, 20.00535, 20.00536, 20.00534, 20.0054, 
    20.00536, 20.00531, 20.00532, 20.00532, 20.00531, 20.00534, 20.00533, 
    20.00536, 20.00535, 20.00537, 20.00536, 20.00536, 20.00535, 20.00535, 
    20.00533, 20.00532, 20.00531, 20.00532, 20.00533, 20.00534, 20.00536, 
    20.00535, 20.00537, 20.00533, 20.00535, 20.00534, 20.00536, 20.00533, 
    20.00535, 20.00532, 20.00533, 20.00533, 20.00535, 20.00535, 20.00536, 
    20.00535, 20.00534, 20.00534, 20.00533, 20.00533, 20.00532, 20.00532, 
    20.00532, 20.00533, 20.00534, 20.00536, 20.00537, 20.00537, 20.00539, 
    20.00538, 20.0054, 20.00538, 20.00541, 20.00535, 20.00538, 20.00533, 
    20.00534, 20.00535, 20.00537, 20.00536, 20.00537, 20.00534, 20.00533, 
    20.00532, 20.00532, 20.00532, 20.00532, 20.00533, 20.00533, 20.00534, 
    20.00533, 20.00536, 20.00537, 20.0054, 20.00541, 20.00543, 20.00544, 
    20.00544, 20.00544,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.525843, 0.5258434, 0.5258433, 0.5258437, 0.5258435, 0.5258437, 0.5258431, 
    0.5258434, 0.5258432, 0.525843, 0.5258443, 0.5258437, 0.525845, 
    0.5258446, 0.5258456, 0.5258449, 0.5258457, 0.5258456, 0.5258461, 
    0.5258459, 0.5258465, 0.5258461, 0.5258468, 0.5258464, 0.5258465, 
    0.5258461, 0.5258438, 0.5258442, 0.5258438, 0.5258439, 0.5258438, 
    0.5258435, 0.5258433, 0.525843, 0.525843, 0.5258433, 0.5258439, 
    0.5258437, 0.5258442, 0.5258442, 0.5258447, 0.5258445, 0.5258454, 
    0.5258451, 0.5258459, 0.5258457, 0.5258459, 0.5258458, 0.5258459, 
    0.5258456, 0.5258458, 0.5258455, 0.5258445, 0.5258448, 0.5258439, 
    0.5258434, 0.5258431, 0.5258428, 0.5258429, 0.525843, 0.5258433, 
    0.5258436, 0.5258439, 0.525844, 0.5258442, 0.5258446, 0.5258449, 
    0.5258455, 0.5258453, 0.5258455, 0.5258457, 0.525846, 0.5258459, 
    0.5258461, 0.5258455, 0.5258459, 0.5258453, 0.5258455, 0.5258442, 
    0.5258437, 0.5258435, 0.5258433, 0.5258429, 0.5258432, 0.5258431, 
    0.5258434, 0.5258436, 0.5258434, 0.525844, 0.5258438, 0.5258449, 
    0.5258445, 0.5258457, 0.5258454, 0.5258458, 0.5258456, 0.5258459, 
    0.5258456, 0.5258461, 0.5258462, 0.5258461, 0.5258464, 0.5258456, 
    0.5258459, 0.5258434, 0.5258435, 0.5258436, 0.5258433, 0.5258432, 
    0.525843, 0.5258432, 0.5258433, 0.5258436, 0.5258437, 0.5258439, 
    0.5258442, 0.5258445, 0.5258451, 0.5258454, 0.5258456, 0.5258455, 
    0.5258456, 0.5258455, 0.5258454, 0.5258462, 0.5258458, 0.5258464, 
    0.5258464, 0.5258461, 0.5258464, 0.5258435, 0.5258434, 0.5258431, 
    0.5258433, 0.5258429, 0.5258431, 0.5258433, 0.5258438, 0.5258439, 
    0.525844, 0.5258442, 0.5258445, 0.5258449, 0.5258453, 0.5258457, 
    0.5258457, 0.5258457, 0.5258458, 0.5258456, 0.5258458, 0.5258458, 
    0.5258458, 0.5258464, 0.5258462, 0.5258464, 0.5258462, 0.5258434, 
    0.5258436, 0.5258435, 0.5258436, 0.5258436, 0.525844, 0.5258441, 
    0.5258448, 0.5258445, 0.5258449, 0.5258445, 0.5258446, 0.5258449, 
    0.5258445, 0.5258453, 0.5258448, 0.5258458, 0.5258452, 0.5258458, 
    0.5258457, 0.5258459, 0.525846, 0.5258462, 0.5258465, 0.5258465, 
    0.5258468, 0.5258438, 0.525844, 0.5258439, 0.5258442, 0.5258443, 
    0.5258446, 0.5258451, 0.5258449, 0.5258452, 0.5258453, 0.5258448, 
    0.5258451, 0.5258441, 0.5258442, 0.5258442, 0.5258438, 0.5258449, 
    0.5258443, 0.5258454, 0.5258451, 0.525846, 0.5258455, 0.5258464, 
    0.5258468, 0.5258472, 0.5258476, 0.525844, 0.5258439, 0.5258442, 
    0.5258445, 0.5258448, 0.5258451, 0.5258452, 0.5258452, 0.5258454, 
    0.5258455, 0.5258452, 0.5258456, 0.5258443, 0.525845, 0.5258439, 
    0.5258442, 0.5258445, 0.5258443, 0.5258449, 0.525845, 0.5258455, 
    0.5258452, 0.5258467, 0.5258461, 0.5258479, 0.5258474, 0.5258439, 
    0.525844, 0.5258446, 0.5258443, 0.5258451, 0.5258453, 0.5258455, 
    0.5258457, 0.5258457, 0.5258458, 0.5258456, 0.5258458, 0.5258451, 
    0.5258454, 0.5258446, 0.5258448, 0.5258447, 0.5258446, 0.5258449, 
    0.5258452, 0.5258452, 0.5258453, 0.5258457, 0.5258451, 0.5258468, 
    0.5258458, 0.5258442, 0.5258446, 0.5258446, 0.5258445, 0.5258453, 
    0.525845, 0.5258458, 0.5258456, 0.5258459, 0.5258458, 0.5258458, 
    0.5258455, 0.5258454, 0.525845, 0.5258448, 0.5258445, 0.5258446, 
    0.5258448, 0.5258453, 0.5258457, 0.5258456, 0.5258459, 0.5258451, 
    0.5258454, 0.5258453, 0.5258456, 0.5258449, 0.5258455, 0.5258447, 
    0.5258448, 0.525845, 0.5258455, 0.5258456, 0.5258456, 0.5258456, 
    0.5258453, 0.5258452, 0.525845, 0.5258449, 0.5258448, 0.5258446, 
    0.5258448, 0.5258449, 0.5258453, 0.5258456, 0.525846, 0.5258461, 
    0.5258466, 0.5258462, 0.5258468, 0.5258463, 0.5258472, 0.5258456, 
    0.5258463, 0.525845, 0.5258452, 0.5258454, 0.5258459, 0.5258456, 
    0.525846, 0.5258452, 0.5258448, 0.5258447, 0.5258445, 0.5258447, 
    0.5258447, 0.5258449, 0.5258448, 0.5258453, 0.5258451, 0.5258458, 
    0.525846, 0.5258468, 0.5258472, 0.5258477, 0.5258479, 0.5258479, 0.525848 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  2.569961e-21, -7.709882e-21, 0, 7.709882e-21, 1.28498e-20, -2.569961e-21, 
    -1.003089e-36, -5.139921e-21, -5.139921e-21, 0, 1.541976e-20, 
    -1.003089e-36, -1.027984e-20, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -1.003089e-36, 1.027984e-20, -7.709882e-21, 1.003089e-36, -7.709882e-21, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, 1.003089e-36, -1.027984e-20, 1.28498e-20, 2.055969e-20, 
    1.003089e-36, -7.709882e-21, -2.569961e-21, -5.139921e-21, -1.798972e-20, 
    -1.003089e-36, -1.003089e-36, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    -2.569961e-21, -1.027984e-20, 1.28498e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -2.569961e-21, 1.027984e-20, -1.027984e-20, -1.541976e-20, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, 7.709882e-21, 1.027984e-20, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -1.28498e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    1.28498e-20, -7.709882e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, 2.569961e-21, -1.28498e-20, -7.709882e-21, -2.569961e-21, 
    -1.541976e-20, 1.28498e-20, -7.709882e-21, 1.003089e-36, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 2.312965e-20, -7.709882e-21, -1.28498e-20, 
    -1.28498e-20, 5.139921e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 1.003089e-36, -1.798972e-20, -1.027984e-20, 2.055969e-20, 
    -1.28498e-20, 7.709882e-21, -5.139921e-21, -1.541976e-20, 0, 
    -2.826957e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 1.027984e-20, 7.709882e-21, -2.312965e-20, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    2.055969e-20, 7.709882e-21, 5.139921e-21, -1.003089e-36, 0, 
    -5.139921e-21, -1.027984e-20, 2.569961e-21, 1.027984e-20, 1.798972e-20, 
    1.027984e-20, 1.541976e-20, 1.027984e-20, -1.798972e-20, 1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, -1.28498e-20, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, -7.709882e-21, 1.003089e-36, 
    -5.139921e-21, 7.709882e-21, 1.027984e-20, 1.28498e-20, 0, -1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, 
    7.709882e-21, 1.027984e-20, 5.139921e-21, 2.826957e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 1.027984e-20, -1.28498e-20, 1.027984e-20, 
    1.798972e-20, 2.569961e-21, -5.139921e-21, -1.541976e-20, 1.027984e-20, 
    -2.569961e-21, -7.709882e-21, -1.798972e-20, 7.709882e-21, -1.541976e-20, 
    -1.28498e-20, -7.709882e-21, -5.139921e-21, 1.541976e-20, -2.569961e-21, 
    -7.709882e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, 0, -1.027984e-20, -7.709882e-21, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, 5.139921e-21, 2.569961e-21, 
    1.28498e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 2.569961e-21, 
    -1.798972e-20, -7.709882e-21, 1.027984e-20, 7.709882e-21, -1.003089e-36, 
    0, 1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    1.027984e-20, 7.709882e-21, -5.139921e-21, -1.798972e-20, -7.709882e-21, 
    -5.139921e-21, -1.027984e-20, -1.541976e-20, 5.139921e-21, -7.709882e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 1.798972e-20, -2.055969e-20, 
    7.709882e-21, 1.027984e-20, 1.28498e-20, -1.003089e-36, 5.139921e-21, 
    -2.569961e-21, 1.541976e-20, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -1.798972e-20, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, -1.003089e-36, 7.709882e-21, 1.027984e-20, -7.709882e-21, 
    -2.569961e-21, 1.28498e-20, -5.139921e-21, -1.28498e-20, 7.709882e-21, 0, 
    -7.709882e-21, 1.003089e-36, -1.541976e-20, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 1.798972e-20, 0, -2.569961e-21, 2.569961e-21, 
    1.027984e-20, -1.28498e-20, 7.709882e-21, 7.709882e-21, -7.709882e-21, 
    -5.139921e-21, -7.709882e-21, -1.28498e-20, -1.003089e-36, -1.027984e-20, 
    1.027984e-20, -1.003089e-36, -1.798972e-20, -5.139921e-21, -1.541976e-20, 
    -2.569961e-21, -5.139921e-21, -1.798972e-20, 1.003089e-36, 1.027984e-20, 
    1.027984e-20, -1.003089e-36, 1.541976e-20, 1.798972e-20, -1.28498e-20, 
    -2.569961e-21, 5.139921e-21, -1.541976e-20, -1.003089e-36, -1.28498e-20, 
    1.28498e-20, -7.709882e-21, 0, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    -1.027984e-20, 2.569961e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -1.28498e-20, 1.003089e-36, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -7.709882e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, -1.28498e-20, 
    3.854941e-20, -1.027984e-20, 2.312965e-20, 5.139921e-21, -1.28498e-20, 
    1.027984e-20, -1.003089e-36, 1.798972e-20, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -2.006177e-36,
  -7.709882e-21, -7.709882e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, 
    -1.541976e-20, 7.709882e-21, -5.139921e-21, 1.003089e-36, -1.541976e-20, 
    -1.003089e-36, -7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, 1.027984e-20, 0, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -1.027984e-20, 1.28498e-20, -1.28498e-20, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -1.28498e-20, 2.569961e-21, 1.027984e-20, 
    1.28498e-20, -2.569961e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -2.569961e-21, 0, 1.003089e-36, 
    5.139921e-21, -2.569961e-21, -1.003089e-36, 0, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, 0, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 0, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, -1.28498e-20, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    7.709882e-21, 1.027984e-20, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, -1.798972e-20, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 1.28498e-20, 1.798972e-20, 
    5.139921e-21, 1.003089e-36, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, -1.541976e-20, -7.709882e-21, -1.003089e-36, -2.569961e-21, 
    -1.027984e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 1.003089e-36, 
    7.709882e-21, -1.798972e-20, -7.709882e-21, -1.28498e-20, 0, 
    -1.541976e-20, 0, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, 0, -2.569961e-21, 1.28498e-20, 0, 
    7.709882e-21, -2.569961e-21, 1.003089e-36, 1.003089e-36, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -1.003089e-36, 1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 2.055969e-20, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 0, 2.569961e-21, -1.003089e-36, 1.541976e-20, 
    -1.003089e-36, 2.569961e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -1.541976e-20, -1.003089e-36, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 1.027984e-20, -1.798972e-20, 2.569961e-21, 1.027984e-20, 
    -1.28498e-20, 2.569961e-21, 0, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 0, -1.027984e-20, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, 0, 5.139921e-21, -1.28498e-20, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, -1.28498e-20, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, 0, -1.027984e-20, 
    1.28498e-20, -2.569961e-21, -2.569961e-21, -2.569961e-21, 0, 0, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -7.709882e-21, -7.709882e-21, 1.541976e-20, 
    7.709882e-21, -1.003089e-36, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -1.28498e-20, 7.709882e-21, -1.28498e-20, 
    -7.709882e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -1.798972e-20, 1.027984e-20, -5.139921e-21, -1.003089e-36, 1.027984e-20, 
    5.139921e-21, 2.569961e-21, -1.28498e-20, 1.027984e-20, -2.569961e-21, 
    7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 0, 
    -1.027984e-20, -5.139921e-21, -1.798972e-20, -2.569961e-21, 7.709882e-21, 
    1.28498e-20, -5.139921e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, 0, -7.709882e-21, 1.003089e-36, 
    -2.569961e-21, 2.569961e-21, 0, -1.027984e-20, -2.569961e-21, 0, 
    -7.709882e-21, 0, -7.709882e-21, 5.139921e-21, 2.569961e-21, 1.28498e-20, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.541976e-20, -2.569961e-21, 
    1.027984e-20, 1.28498e-20, 1.003089e-36, 5.139921e-21, 0, -2.569961e-21, 
    1.003089e-36, -1.027984e-20, -2.569961e-21, 0, -1.003089e-36, 
    -1.003089e-36, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    1.798972e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, -1.798972e-20, -5.139921e-21, 1.027984e-20, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, 0, -7.709882e-21, 
    -2.569961e-21, 0, -1.28498e-20, 7.709882e-21, 1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 0, -1.027984e-20, 0, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 0, -2.569961e-21, 5.139921e-21, -2.569961e-21,
  1.28498e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 2.569961e-21, 
    -7.709882e-21, -1.003089e-36, -7.709882e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.003089e-36, 0, 0, 1.027984e-20, 7.709882e-21, 
    1.541976e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    1.027984e-20, -1.027984e-20, 5.139921e-21, -1.28498e-20, 0, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 1.003089e-36, 2.569961e-21, 
    -1.003089e-36, -1.541976e-20, 5.139921e-21, 1.027984e-20, 0, 
    2.569961e-21, 7.709882e-21, -1.541976e-20, 2.569961e-21, -1.027984e-20, 
    -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    1.003089e-36, -2.569961e-21, 0, -2.569961e-21, 1.027984e-20, 
    1.798972e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 5.139921e-21, 
    2.569961e-21, -1.027984e-20, -5.139921e-21, 0, -1.28498e-20, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 2.055969e-20, 5.139921e-21, -2.569961e-21, 
    1.798972e-20, 2.569961e-21, -1.28498e-20, 0, -1.28498e-20, 5.139921e-21, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 1.28498e-20, 7.709882e-21, -1.027984e-20, 
    1.003089e-36, -1.027984e-20, 5.139921e-21, 1.28498e-20, 0, 2.826957e-20, 
    -1.003089e-36, -2.569961e-21, -1.28498e-20, -1.027984e-20, 0, 
    -5.139921e-21, 2.569961e-21, 1.003089e-36, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, -2.569961e-21, -7.709882e-21, 1.003089e-36, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, -1.003089e-36, 
    -2.569961e-21, 5.139921e-21, 1.003089e-36, 2.569961e-21, -1.027984e-20, 
    1.798972e-20, -5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -1.798972e-20, -2.569961e-21, 0, 2.569961e-21, 1.28498e-20, 5.139921e-21, 
    -2.569961e-21, -5.139921e-21, 0, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, -1.28498e-20, 1.027984e-20, 
    5.139921e-21, 0, 1.541976e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    1.798972e-20, 2.569961e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, 1.027984e-20, -7.709882e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 0, 
    -1.003089e-36, 2.569961e-21, 7.709882e-21, 1.027984e-20, 0, -1.28498e-20, 
    0, 2.569961e-21, 2.569961e-21, -5.139921e-21, -1.027984e-20, 
    1.798972e-20, 5.139921e-21, 7.709882e-21, -7.709882e-21, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, -2.569961e-21, -7.709882e-21, 
    -1.798972e-20, 7.709882e-21, -7.709882e-21, 1.003089e-36, 5.139921e-21, 
    -1.28498e-20, 5.139921e-21, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    -7.709882e-21, 0, 0, 5.139921e-21, -1.28498e-20, -1.027984e-20, 
    -1.541976e-20, -7.709882e-21, 1.28498e-20, 0, -5.139921e-21, 1.28498e-20, 
    0, -7.709882e-21, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    1.28498e-20, -1.541976e-20, 1.027984e-20, 7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, 0, -1.027984e-20, 2.569961e-21, 0, 
    -2.569961e-21, 2.569961e-21, -1.798972e-20, 1.003089e-36, 0, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 1.28498e-20, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, 0, -1.003089e-36, 
    7.709882e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    7.709882e-21, 0, -1.28498e-20, 0, 2.569961e-21, 5.139921e-21, 
    1.003089e-36, 0, -1.003089e-36, 1.003089e-36, -2.569961e-21, 1.28498e-20, 
    2.569961e-21, 0, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, 0, -1.003089e-36, -1.28498e-20, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 5.139921e-21, 0, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 0, -2.569961e-21, 
    -1.541976e-20, -2.312965e-20, 1.28498e-20, 7.709882e-21, 1.027984e-20, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, -1.003089e-36, -2.569961e-21, 
    7.709882e-21, 1.28498e-20, 0, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    1.003089e-36, 7.709882e-21, 7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, -1.541976e-20, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 
    -1.027984e-20, 5.139921e-21, 1.027984e-20, -1.003089e-36, -7.709882e-21, 
    7.709882e-21, 1.28498e-20, -5.139921e-21, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, 0, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, -1.541976e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 0, -1.027984e-20,
  1.027984e-20, -1.027984e-20, 2.569961e-21, 0, 2.569961e-21, 2.055969e-20, 
    5.139921e-21, 0, -1.027984e-20, 7.709882e-21, -5.139921e-21, 
    -1.003089e-36, 2.569961e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -2.569961e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 0, -2.055969e-20, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, 7.709882e-21, -2.569961e-20, 1.798972e-20, 
    1.003089e-36, -5.139921e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 1.28498e-20, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -1.027984e-20, 1.027984e-20, 7.709882e-21, 
    -2.569961e-21, 1.027984e-20, 0, -2.569961e-21, -1.28498e-20, 0, 
    -5.139921e-21, 1.28498e-20, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -1.28498e-20, 0, -1.027984e-20, 1.027984e-20, 1.28498e-20, 
    -1.027984e-20, 7.709882e-21, 1.027984e-20, 7.709882e-21, 1.28498e-20, 
    -1.027984e-20, -1.003089e-36, -5.139921e-21, -1.541976e-20, -1.28498e-20, 
    -2.055969e-20, -5.139921e-21, 2.569961e-21, -5.139921e-21, -1.003089e-36, 
    5.139921e-21, 7.709882e-21, -1.28498e-20, 5.139921e-21, 1.28498e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, -1.798972e-20, -1.28498e-20, 
    1.027984e-20, -2.569961e-21, -7.709882e-21, -2.569961e-21, -1.003089e-36, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, 0, -2.055969e-20, 
    1.541976e-20, -1.003089e-36, 1.798972e-20, 2.569961e-21, -5.139921e-21, 
    -1.003089e-36, -1.027984e-20, -5.139921e-21, 1.027984e-20, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    1.027984e-20, -5.139921e-21, -2.312965e-20, 2.569961e-21, 1.003089e-36, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -1.28498e-20, 2.055969e-20, 1.541976e-20, -1.798972e-20, 1.027984e-20, 
    1.541976e-20, -1.003089e-36, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    7.709882e-21, -1.28498e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, 
    0, -7.709882e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 7.709882e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -1.541976e-20, 2.569961e-21, 1.027984e-20, -2.055969e-20, -7.709882e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 1.027984e-20, 
    1.003089e-36, 1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -1.28498e-20, 0, -1.003089e-36, -1.003089e-36, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 1.003089e-36, -7.709882e-21, -1.541976e-20, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, -1.28498e-20, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, -1.798972e-20, 0, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    0, 7.709882e-21, 2.569961e-21, -1.28498e-20, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, -7.709882e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, -1.541976e-20, 
    7.709882e-21, -1.027984e-20, -1.28498e-20, 1.027984e-20, -2.569961e-21, 
    -1.541976e-20, -1.28498e-20, 2.569961e-21, -5.139921e-21, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, -1.003089e-36, 1.027984e-20, 
    -7.709882e-21, 7.709882e-21, -1.28498e-20, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, -2.312965e-20, 2.569961e-21, 2.569961e-21, 1.28498e-20, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, 1.003089e-36, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 1.003089e-36, -1.28498e-20, -1.027984e-20, -1.28498e-20, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    1.027984e-20, -7.709882e-21, -2.569961e-21, 1.027984e-20, -2.826957e-20, 
    -7.709882e-21, -7.709882e-21, -1.28498e-20, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 7.709882e-21, 1.541976e-20, 5.139921e-21, 
    1.003089e-36, 7.709882e-21, -5.139921e-21, 0, -1.798972e-20, 
    -1.003089e-36, 5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 0, -1.003089e-36, 1.28498e-20, 7.709882e-21, 
    -2.055969e-20, -1.003089e-36, 7.709882e-21, -7.709882e-21, 7.709882e-21, 
    -1.027984e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 1.541976e-20, 5.139921e-21, 1.28498e-20, 0, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 0,
  -5.139921e-21, 5.139921e-21, -5.139921e-21, 0, 2.569961e-21, -1.798972e-20, 
    -1.003089e-36, 1.003089e-36, 1.027984e-20, 1.003089e-36, 1.28498e-20, 
    5.139921e-21, 2.569961e-21, -7.709882e-21, -1.003089e-36, 1.541976e-20, 
    2.569961e-21, 1.027984e-20, -1.28498e-20, -2.312965e-20, 1.28498e-20, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, 1.541976e-20, -2.569961e-21, 
    2.312965e-20, 1.027984e-20, -1.541976e-20, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.027984e-20, 1.541976e-20, 7.709882e-21, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, 1.027984e-20, 7.709882e-21, 1.28498e-20, 
    5.139921e-21, 2.569961e-21, -2.569961e-20, -7.709882e-21, -3.083953e-20, 
    -1.003089e-36, 2.569961e-21, 5.139921e-21, 0, 1.28498e-20, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, 2.055969e-20, 
    -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, -1.003089e-36, 
    -1.28498e-20, 5.139921e-21, 2.569961e-21, -1.003089e-36, -1.027984e-20, 
    1.798972e-20, -1.027984e-20, -5.139921e-21, -5.139921e-21, 1.28498e-20, 
    1.027984e-20, -7.709882e-21, 2.569961e-21, -1.28498e-20, -1.027984e-20, 
    -1.003089e-36, -1.027984e-20, 1.798972e-20, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, 2.055969e-20, 2.569961e-21, -2.569961e-21, -1.798972e-20, 
    -7.709882e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, -1.003089e-36, 1.28498e-20, -5.139921e-21, -5.139921e-21, 
    -1.28498e-20, 1.28498e-20, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, 1.027984e-20, 1.28498e-20, 1.027984e-20, 1.003089e-36, 
    -1.027984e-20, -1.541976e-20, -1.003089e-36, -5.139921e-21, 
    -7.709882e-21, 5.139921e-21, 2.055969e-20, -1.798972e-20, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 1.28498e-20, 7.709882e-21, 0, -7.709882e-21, 
    7.709882e-21, -1.28498e-20, -1.027984e-20, 0, 2.569961e-21, 
    -2.569961e-21, 1.28498e-20, -2.569961e-21, -5.139921e-21, -1.027984e-20, 
    7.709882e-21, 1.28498e-20, 0, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -3.009266e-36, -5.139921e-21, 1.003089e-36, -7.709882e-21, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, 2.312965e-20, 
    -1.541976e-20, -2.055969e-20, 1.027984e-20, -1.798972e-20, -2.569961e-21, 
    -2.312965e-20, -5.139921e-21, -7.709882e-21, 1.003089e-36, 2.569961e-21, 
    -5.139921e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, -1.28498e-20, 
    -2.055969e-20, 2.055969e-20, 1.798972e-20, 5.139921e-21, 7.709882e-21, 
    7.709882e-21, -5.139921e-21, 7.709882e-21, 1.28498e-20, -1.798972e-20, 
    2.312965e-20, 1.541976e-20, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, 7.709882e-21, 2.055969e-20, 
    -1.027984e-20, 1.28498e-20, 7.709882e-21, 5.139921e-21, 1.798972e-20, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, 1.027984e-20, 2.569961e-21, -2.569961e-21, 1.28498e-20, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, -1.027984e-20, 2.569961e-21, 
    -2.826957e-20, -1.798972e-20, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -1.28498e-20, 7.709882e-21, 7.709882e-21, 1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, 1.28498e-20, 5.139921e-21, 1.541976e-20, 1.027984e-20, 
    -1.541976e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 1.798972e-20, 
    2.055969e-20, -7.709882e-21, 2.569961e-21, 0, 1.541976e-20, 
    -1.003089e-36, -2.569961e-20, -1.541976e-20, 7.709882e-21, -1.541976e-20, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, 7.709882e-21, 
    1.003089e-36, -1.541976e-20, 1.28498e-20, 7.709882e-21, 1.798972e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, 
    0, 7.709882e-21, 1.027984e-20, -1.541976e-20, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-20, 1.28498e-20, -1.28498e-20, -1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 2.312965e-20, -5.139921e-21, -7.709882e-21, 
    1.027984e-20, 1.003089e-36, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 1.28498e-20, -5.139921e-21, -1.003089e-36, -7.709882e-21, 
    -5.139921e-21, 1.798972e-20, 1.003089e-36, -7.709882e-21, -1.28498e-20, 
    7.709882e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, -1.28498e-20, 
    1.027984e-20, -7.709882e-21, -5.139921e-21, 1.541976e-20, 2.055969e-20, 
    7.709882e-21, 2.569961e-21, 2.055969e-20, 1.003089e-36, 1.027984e-20, 
    1.28498e-20, -1.003089e-36, -2.569961e-21, -3.083953e-20, -1.003089e-36, 
    1.798972e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 
    -7.709882e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, -1.798972e-20, 1.541976e-20, -7.709882e-21, -1.003089e-36, 
    1.798972e-20, -1.28498e-20, -1.798972e-20, 1.798972e-20,
  6.259692e-29, 6.259697e-29, 6.259697e-29, 6.2597e-29, 6.259698e-29, 
    6.2597e-29, 6.259694e-29, 6.259697e-29, 6.259695e-29, 6.259693e-29, 
    6.259707e-29, 6.2597e-29, 6.259715e-29, 6.25971e-29, 6.259721e-29, 
    6.259714e-29, 6.259723e-29, 6.259721e-29, 6.259727e-29, 6.259725e-29, 
    6.259732e-29, 6.259727e-29, 6.259735e-29, 6.259731e-29, 6.259732e-29, 
    6.259727e-29, 6.259701e-29, 6.259706e-29, 6.259701e-29, 6.259702e-29, 
    6.259702e-29, 6.259698e-29, 6.259696e-29, 6.259692e-29, 6.259693e-29, 
    6.259696e-29, 6.259703e-29, 6.2597e-29, 6.259706e-29, 6.259706e-29, 
    6.259712e-29, 6.259709e-29, 6.259719e-29, 6.259716e-29, 6.259725e-29, 
    6.259723e-29, 6.259725e-29, 6.259724e-29, 6.259725e-29, 6.259722e-29, 
    6.259723e-29, 6.259721e-29, 6.25971e-29, 6.259713e-29, 6.259703e-29, 
    6.259698e-29, 6.259694e-29, 6.259691e-29, 6.259691e-29, 6.259692e-29, 
    6.259696e-29, 6.2597e-29, 6.259702e-29, 6.259704e-29, 6.259706e-29, 
    6.259711e-29, 6.259714e-29, 6.25972e-29, 6.259719e-29, 6.259721e-29, 
    6.259723e-29, 6.259726e-29, 6.259726e-29, 6.259727e-29, 6.259721e-29, 
    6.259725e-29, 6.259718e-29, 6.25972e-29, 6.259706e-29, 6.259701e-29, 
    6.259698e-29, 6.259697e-29, 6.259692e-29, 6.259695e-29, 6.259694e-29, 
    6.259697e-29, 6.259699e-29, 6.259698e-29, 6.259704e-29, 6.259701e-29, 
    6.259714e-29, 6.259709e-29, 6.259723e-29, 6.259719e-29, 6.259723e-29, 
    6.259721e-29, 6.259725e-29, 6.259722e-29, 6.259727e-29, 6.259729e-29, 
    6.259728e-29, 6.259731e-29, 6.259721e-29, 6.259725e-29, 6.259698e-29, 
    6.259698e-29, 6.259699e-29, 6.259695e-29, 6.259695e-29, 6.259692e-29, 
    6.259695e-29, 6.259696e-29, 6.259699e-29, 6.259701e-29, 6.259702e-29, 
    6.259706e-29, 6.25971e-29, 6.259715e-29, 6.259719e-29, 6.259722e-29, 
    6.259721e-29, 6.259722e-29, 6.25972e-29, 6.259719e-29, 6.259728e-29, 
    6.259723e-29, 6.25973e-29, 6.25973e-29, 6.259727e-29, 6.25973e-29, 
    6.259698e-29, 6.259697e-29, 6.259694e-29, 6.259697e-29, 6.259692e-29, 
    6.259694e-29, 6.259696e-29, 6.259701e-29, 6.259703e-29, 6.259704e-29, 
    6.259706e-29, 6.259709e-29, 6.259714e-29, 6.259719e-29, 6.259723e-29, 
    6.259723e-29, 6.259723e-29, 6.259724e-29, 6.259721e-29, 6.259724e-29, 
    6.259724e-29, 6.259723e-29, 6.25973e-29, 6.259728e-29, 6.25973e-29, 
    6.259729e-29, 6.259697e-29, 6.259699e-29, 6.259698e-29, 6.2597e-29, 
    6.259698e-29, 6.259704e-29, 6.259705e-29, 6.259712e-29, 6.259709e-29, 
    6.259713e-29, 6.25971e-29, 6.25971e-29, 6.259714e-29, 6.25971e-29, 
    6.259718e-29, 6.259713e-29, 6.259724e-29, 6.259718e-29, 6.259724e-29, 
    6.259723e-29, 6.259725e-29, 6.259727e-29, 6.259729e-29, 6.259733e-29, 
    6.259732e-29, 6.259735e-29, 6.259701e-29, 6.259703e-29, 6.259703e-29, 
    6.259705e-29, 6.259707e-29, 6.25971e-29, 6.259716e-29, 6.259713e-29, 
    6.259717e-29, 6.259718e-29, 6.259712e-29, 6.259716e-29, 6.259704e-29, 
    6.259706e-29, 6.259706e-29, 6.259701e-29, 6.259714e-29, 6.259707e-29, 
    6.259719e-29, 6.259716e-29, 6.259726e-29, 6.259721e-29, 6.259731e-29, 
    6.259735e-29, 6.259739e-29, 6.259744e-29, 6.259704e-29, 6.259703e-29, 
    6.259706e-29, 6.259709e-29, 6.259712e-29, 6.259716e-29, 6.259716e-29, 
    6.259718e-29, 6.259719e-29, 6.259721e-29, 6.259718e-29, 6.259722e-29, 
    6.259707e-29, 6.259715e-29, 6.259703e-29, 6.259706e-29, 6.259709e-29, 
    6.259707e-29, 6.259713e-29, 6.259715e-29, 6.25972e-29, 6.259717e-29, 
    6.259735e-29, 6.259727e-29, 6.259748e-29, 6.259742e-29, 6.259703e-29, 
    6.259704e-29, 6.259711e-29, 6.259708e-29, 6.259716e-29, 6.259719e-29, 
    6.259721e-29, 6.259723e-29, 6.259723e-29, 6.259724e-29, 6.259722e-29, 
    6.259724e-29, 6.259716e-29, 6.259719e-29, 6.25971e-29, 6.259712e-29, 
    6.259712e-29, 6.25971e-29, 6.259714e-29, 6.259718e-29, 6.259718e-29, 
    6.259719e-29, 6.259723e-29, 6.259716e-29, 6.259735e-29, 6.259724e-29, 
    6.259706e-29, 6.25971e-29, 6.25971e-29, 6.259709e-29, 6.259718e-29, 
    6.259715e-29, 6.259724e-29, 6.259722e-29, 6.259726e-29, 6.259724e-29, 
    6.259724e-29, 6.259721e-29, 6.259719e-29, 6.259715e-29, 6.259712e-29, 
    6.259709e-29, 6.25971e-29, 6.259713e-29, 6.259718e-29, 6.259723e-29, 
    6.259722e-29, 6.259726e-29, 6.259716e-29, 6.25972e-29, 6.259718e-29, 
    6.259723e-29, 6.259713e-29, 6.259721e-29, 6.259712e-29, 6.259712e-29, 
    6.259715e-29, 6.25972e-29, 6.259721e-29, 6.259723e-29, 6.259722e-29, 
    6.259718e-29, 6.259718e-29, 6.259715e-29, 6.259714e-29, 6.259712e-29, 
    6.25971e-29, 6.259712e-29, 6.259713e-29, 6.259718e-29, 6.259722e-29, 
    6.259727e-29, 6.259727e-29, 6.259733e-29, 6.259729e-29, 6.259735e-29, 
    6.25973e-29, 6.259739e-29, 6.259721e-29, 6.259729e-29, 6.259715e-29, 
    6.259716e-29, 6.259719e-29, 6.259726e-29, 6.259723e-29, 6.259726e-29, 
    6.259718e-29, 6.259713e-29, 6.259712e-29, 6.259709e-29, 6.259712e-29, 
    6.259712e-29, 6.259713e-29, 6.259713e-29, 6.259718e-29, 6.259715e-29, 
    6.259724e-29, 6.259726e-29, 6.259735e-29, 6.259739e-29, 6.259745e-29, 
    6.259747e-29, 6.259748e-29, 6.259748e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.631813e-10, 2.639023e-10, 2.637622e-10, 2.643435e-10, 2.640211e-10, 
    2.644017e-10, 2.633275e-10, 2.639308e-10, 2.635457e-10, 2.632463e-10, 
    2.654712e-10, 2.643695e-10, 2.666157e-10, 2.659133e-10, 2.676776e-10, 
    2.665064e-10, 2.679137e-10, 2.676439e-10, 2.684561e-10, 2.682235e-10, 
    2.692618e-10, 2.685635e-10, 2.698001e-10, 2.690952e-10, 2.692054e-10, 
    2.685405e-10, 2.645913e-10, 2.653341e-10, 2.645473e-10, 2.646532e-10, 
    2.646057e-10, 2.640277e-10, 2.637363e-10, 2.631262e-10, 2.63237e-10, 
    2.636851e-10, 2.647009e-10, 2.643562e-10, 2.65225e-10, 2.652054e-10, 
    2.661723e-10, 2.657363e-10, 2.67361e-10, 2.668994e-10, 2.682332e-10, 
    2.678978e-10, 2.682174e-10, 2.681205e-10, 2.682187e-10, 2.677268e-10, 
    2.679375e-10, 2.675047e-10, 2.65818e-10, 2.663137e-10, 2.648347e-10, 
    2.639449e-10, 2.633539e-10, 2.629345e-10, 2.629938e-10, 2.631068e-10, 
    2.636877e-10, 2.642339e-10, 2.646501e-10, 2.649284e-10, 2.652026e-10, 
    2.660321e-10, 2.664713e-10, 2.674543e-10, 2.67277e-10, 2.675774e-10, 
    2.678645e-10, 2.683462e-10, 2.682669e-10, 2.684791e-10, 2.675695e-10, 
    2.68174e-10, 2.67176e-10, 2.67449e-10, 2.652767e-10, 2.644492e-10, 
    2.64097e-10, 2.637891e-10, 2.630394e-10, 2.635571e-10, 2.63353e-10, 
    2.638386e-10, 2.641471e-10, 2.639945e-10, 2.64936e-10, 2.6457e-10, 
    2.664973e-10, 2.656673e-10, 2.67831e-10, 2.673134e-10, 2.67955e-10, 
    2.676276e-10, 2.681885e-10, 2.676838e-10, 2.685581e-10, 2.687484e-10, 
    2.686184e-10, 2.691181e-10, 2.676558e-10, 2.682174e-10, 2.639902e-10, 
    2.640151e-10, 2.641311e-10, 2.636214e-10, 2.635902e-10, 2.631232e-10, 
    2.635388e-10, 2.637157e-10, 2.64165e-10, 2.644306e-10, 2.646831e-10, 
    2.652382e-10, 2.65858e-10, 2.667245e-10, 2.67347e-10, 2.677641e-10, 
    2.675083e-10, 2.677341e-10, 2.674817e-10, 2.673634e-10, 2.686771e-10, 
    2.679395e-10, 2.690462e-10, 2.68985e-10, 2.684842e-10, 2.689919e-10, 
    2.640326e-10, 2.638894e-10, 2.633922e-10, 2.637813e-10, 2.630723e-10, 
    2.634692e-10, 2.636973e-10, 2.645776e-10, 2.64771e-10, 2.649503e-10, 
    2.653044e-10, 2.657587e-10, 2.665554e-10, 2.672485e-10, 2.678812e-10, 
    2.678348e-10, 2.678511e-10, 2.679924e-10, 2.676424e-10, 2.680498e-10, 
    2.681182e-10, 2.679394e-10, 2.689768e-10, 2.686805e-10, 2.689837e-10, 
    2.687908e-10, 2.63936e-10, 2.641769e-10, 2.640467e-10, 2.642915e-10, 
    2.64119e-10, 2.648857e-10, 2.651156e-10, 2.661908e-10, 2.657497e-10, 
    2.664519e-10, 2.658211e-10, 2.659328e-10, 2.664746e-10, 2.658552e-10, 
    2.672102e-10, 2.662915e-10, 2.679979e-10, 2.670805e-10, 2.680554e-10, 
    2.678784e-10, 2.681714e-10, 2.684337e-10, 2.687638e-10, 2.693725e-10, 
    2.692316e-10, 2.697407e-10, 2.64536e-10, 2.648484e-10, 2.64821e-10, 
    2.651478e-10, 2.653896e-10, 2.659135e-10, 2.667536e-10, 2.664378e-10, 
    2.670176e-10, 2.67134e-10, 2.66253e-10, 2.667939e-10, 2.650575e-10, 
    2.65338e-10, 2.65171e-10, 2.645606e-10, 2.665104e-10, 2.655099e-10, 
    2.673572e-10, 2.668154e-10, 2.683963e-10, 2.676102e-10, 2.69154e-10, 
    2.698135e-10, 2.704344e-10, 2.711594e-10, 2.650189e-10, 2.648067e-10, 
    2.651868e-10, 2.657124e-10, 2.662002e-10, 2.668485e-10, 2.669148e-10, 
    2.670362e-10, 2.673508e-10, 2.676152e-10, 2.670746e-10, 2.676814e-10, 
    2.654029e-10, 2.665973e-10, 2.647264e-10, 2.652898e-10, 2.656814e-10, 
    2.655097e-10, 2.664017e-10, 2.666118e-10, 2.674656e-10, 2.670243e-10, 
    2.696507e-10, 2.68489e-10, 2.717116e-10, 2.708114e-10, 2.647325e-10, 
    2.650182e-10, 2.660123e-10, 2.655394e-10, 2.668918e-10, 2.672245e-10, 
    2.674951e-10, 2.678407e-10, 2.678781e-10, 2.680829e-10, 2.677473e-10, 
    2.680697e-10, 2.668498e-10, 2.673951e-10, 2.658987e-10, 2.66263e-10, 
    2.660955e-10, 2.659116e-10, 2.664789e-10, 2.670831e-10, 2.670961e-10, 
    2.672897e-10, 2.678352e-10, 2.668973e-10, 2.698003e-10, 2.680077e-10, 
    2.653298e-10, 2.658798e-10, 2.659584e-10, 2.657454e-10, 2.671912e-10, 
    2.666674e-10, 2.680779e-10, 2.676968e-10, 2.683213e-10, 2.68011e-10, 
    2.679653e-10, 2.675667e-10, 2.673185e-10, 2.666914e-10, 2.66181e-10, 
    2.657763e-10, 2.658704e-10, 2.66315e-10, 2.6712e-10, 2.678814e-10, 
    2.677147e-10, 2.682738e-10, 2.667938e-10, 2.674144e-10, 2.671745e-10, 
    2.678e-10, 2.664294e-10, 2.675962e-10, 2.661309e-10, 2.662595e-10, 
    2.66657e-10, 2.674564e-10, 2.676334e-10, 2.678222e-10, 2.677057e-10, 
    2.671405e-10, 2.670479e-10, 2.666474e-10, 2.665367e-10, 2.662315e-10, 
    2.659787e-10, 2.662096e-10, 2.664521e-10, 2.671408e-10, 2.677612e-10, 
    2.684374e-10, 2.686029e-10, 2.693925e-10, 2.687497e-10, 2.698103e-10, 
    2.689084e-10, 2.704696e-10, 2.67664e-10, 2.68882e-10, 2.666751e-10, 
    2.66913e-10, 2.673431e-10, 2.683294e-10, 2.677971e-10, 2.684197e-10, 
    2.670443e-10, 2.663303e-10, 2.661456e-10, 2.658009e-10, 2.661535e-10, 
    2.661248e-10, 2.664622e-10, 2.663538e-10, 2.671636e-10, 2.667287e-10, 
    2.679642e-10, 2.684148e-10, 2.696873e-10, 2.70467e-10, 2.712606e-10, 
    2.716109e-10, 2.717175e-10, 2.717621e-10 ;

 SOIL2N_TO_SOIL3N =
  1.879866e-11, 1.885016e-11, 1.884016e-11, 1.888168e-11, 1.885865e-11, 
    1.888584e-11, 1.880911e-11, 1.88522e-11, 1.88247e-11, 1.88033e-11, 
    1.896223e-11, 1.888353e-11, 1.904398e-11, 1.899381e-11, 1.911983e-11, 
    1.903617e-11, 1.913669e-11, 1.911742e-11, 1.917544e-11, 1.915882e-11, 
    1.923299e-11, 1.918311e-11, 1.927144e-11, 1.922108e-11, 1.922896e-11, 
    1.918146e-11, 1.889938e-11, 1.895243e-11, 1.889624e-11, 1.89038e-11, 
    1.890041e-11, 1.885912e-11, 1.883831e-11, 1.879473e-11, 1.880265e-11, 
    1.883465e-11, 1.89072e-11, 1.888258e-11, 1.894464e-11, 1.894324e-11, 
    1.90123e-11, 1.898117e-11, 1.909721e-11, 1.906424e-11, 1.915951e-11, 
    1.913556e-11, 1.915839e-11, 1.915147e-11, 1.915848e-11, 1.912334e-11, 
    1.91384e-11, 1.910748e-11, 1.8987e-11, 1.902241e-11, 1.891677e-11, 
    1.885321e-11, 1.8811e-11, 1.878103e-11, 1.878527e-11, 1.879334e-11, 
    1.883484e-11, 1.887385e-11, 1.890357e-11, 1.892345e-11, 1.894304e-11, 
    1.900229e-11, 1.903367e-11, 1.910387e-11, 1.909121e-11, 1.911267e-11, 
    1.913317e-11, 1.916758e-11, 1.916192e-11, 1.917708e-11, 1.911211e-11, 
    1.915529e-11, 1.9084e-11, 1.91035e-11, 1.894834e-11, 1.888923e-11, 
    1.886408e-11, 1.884208e-11, 1.878853e-11, 1.882551e-11, 1.881093e-11, 
    1.884561e-11, 1.886765e-11, 1.885675e-11, 1.8924e-11, 1.889786e-11, 
    1.903552e-11, 1.897624e-11, 1.913078e-11, 1.909381e-11, 1.913964e-11, 
    1.911626e-11, 1.915632e-11, 1.912027e-11, 1.918272e-11, 1.919632e-11, 
    1.918703e-11, 1.922272e-11, 1.911827e-11, 1.915838e-11, 1.885645e-11, 
    1.885822e-11, 1.88665e-11, 1.88301e-11, 1.882787e-11, 1.879451e-11, 
    1.88242e-11, 1.883684e-11, 1.886893e-11, 1.88879e-11, 1.890594e-11, 
    1.894559e-11, 1.898986e-11, 1.905175e-11, 1.909621e-11, 1.9126e-11, 
    1.910774e-11, 1.912386e-11, 1.910583e-11, 1.909739e-11, 1.919122e-11, 
    1.913854e-11, 1.921759e-11, 1.921322e-11, 1.917744e-11, 1.921371e-11, 
    1.885947e-11, 1.884925e-11, 1.881373e-11, 1.884152e-11, 1.879088e-11, 
    1.881923e-11, 1.883552e-11, 1.88984e-11, 1.891222e-11, 1.892502e-11, 
    1.895031e-11, 1.898276e-11, 1.903967e-11, 1.908918e-11, 1.913437e-11, 
    1.913106e-11, 1.913222e-11, 1.914231e-11, 1.911732e-11, 1.914642e-11, 
    1.91513e-11, 1.913853e-11, 1.921263e-11, 1.919146e-11, 1.921312e-11, 
    1.919934e-11, 1.885257e-11, 1.886978e-11, 1.886048e-11, 1.887796e-11, 
    1.886564e-11, 1.892041e-11, 1.893683e-11, 1.901363e-11, 1.898212e-11, 
    1.903228e-11, 1.898722e-11, 1.89952e-11, 1.90339e-11, 1.898966e-11, 
    1.908645e-11, 1.902082e-11, 1.91427e-11, 1.907718e-11, 1.914681e-11, 
    1.913417e-11, 1.91551e-11, 1.917384e-11, 1.919741e-11, 1.92409e-11, 
    1.923083e-11, 1.926719e-11, 1.889543e-11, 1.891774e-11, 1.891578e-11, 
    1.893913e-11, 1.89564e-11, 1.899382e-11, 1.905383e-11, 1.903127e-11, 
    1.907269e-11, 1.9081e-11, 1.901808e-11, 1.905671e-11, 1.893268e-11, 
    1.895272e-11, 1.894079e-11, 1.889719e-11, 1.903646e-11, 1.896499e-11, 
    1.909694e-11, 1.905825e-11, 1.917116e-11, 1.911501e-11, 1.922529e-11, 
    1.927239e-11, 1.931674e-11, 1.936853e-11, 1.892992e-11, 1.891476e-11, 
    1.894191e-11, 1.897946e-11, 1.90143e-11, 1.90606e-11, 1.906534e-11, 
    1.907402e-11, 1.909648e-11, 1.911537e-11, 1.907675e-11, 1.91201e-11, 
    1.895735e-11, 1.904266e-11, 1.890903e-11, 1.894927e-11, 1.897725e-11, 
    1.896498e-11, 1.902869e-11, 1.90437e-11, 1.910469e-11, 1.907317e-11, 
    1.926076e-11, 1.917779e-11, 1.940797e-11, 1.934367e-11, 1.890947e-11, 
    1.892987e-11, 1.900088e-11, 1.89671e-11, 1.90637e-11, 1.908747e-11, 
    1.910679e-11, 1.913148e-11, 1.913415e-11, 1.914878e-11, 1.912481e-11, 
    1.914783e-11, 1.90607e-11, 1.909965e-11, 1.899277e-11, 1.901878e-11, 
    1.900682e-11, 1.899369e-11, 1.903421e-11, 1.907736e-11, 1.907829e-11, 
    1.909212e-11, 1.913108e-11, 1.906409e-11, 1.927145e-11, 1.914341e-11, 
    1.895212e-11, 1.899141e-11, 1.899703e-11, 1.898181e-11, 1.908508e-11, 
    1.904767e-11, 1.914842e-11, 1.91212e-11, 1.91658e-11, 1.914364e-11, 
    1.914038e-11, 1.911191e-11, 1.909418e-11, 1.904939e-11, 1.901293e-11, 
    1.898402e-11, 1.899074e-11, 1.90225e-11, 1.908e-11, 1.913439e-11, 
    1.912248e-11, 1.916242e-11, 1.90567e-11, 1.910103e-11, 1.908389e-11, 
    1.912857e-11, 1.903067e-11, 1.911402e-11, 1.900935e-11, 1.901853e-11, 
    1.904693e-11, 1.910403e-11, 1.911667e-11, 1.913016e-11, 1.912184e-11, 
    1.908146e-11, 1.907485e-11, 1.904624e-11, 1.903834e-11, 1.901653e-11, 
    1.899848e-11, 1.901497e-11, 1.903229e-11, 1.908148e-11, 1.91258e-11, 
    1.91741e-11, 1.918593e-11, 1.924232e-11, 1.91964e-11, 1.927217e-11, 
    1.920774e-11, 1.931926e-11, 1.911886e-11, 1.920586e-11, 1.904822e-11, 
    1.906521e-11, 1.909593e-11, 1.916639e-11, 1.912836e-11, 1.917284e-11, 
    1.907459e-11, 1.902359e-11, 1.90104e-11, 1.898578e-11, 1.901096e-11, 
    1.900892e-11, 1.903302e-11, 1.902527e-11, 1.908312e-11, 1.905205e-11, 
    1.91403e-11, 1.917249e-11, 1.926338e-11, 1.931907e-11, 1.937576e-11, 
    1.940078e-11, 1.940839e-11, 1.941157e-11 ;

 SOIL2N_vr =
  1.818739, 1.81874, 1.81874, 1.818741, 1.81874, 1.818741, 1.818739, 1.81874, 
    1.818739, 1.818739, 1.818743, 1.818741, 1.818745, 1.818744, 1.818748, 
    1.818745, 1.818748, 1.818748, 1.818749, 1.818749, 1.818751, 1.818749, 
    1.818752, 1.81875, 1.818751, 1.818749, 1.818741, 1.818743, 1.818741, 
    1.818742, 1.818742, 1.81874, 1.81874, 1.818739, 1.818739, 1.81874, 
    1.818742, 1.818741, 1.818743, 1.818743, 1.818745, 1.818744, 1.818747, 
    1.818746, 1.818749, 1.818748, 1.818749, 1.818748, 1.818749, 1.818748, 
    1.818748, 1.818747, 1.818744, 1.818745, 1.818742, 1.81874, 1.818739, 
    1.818738, 1.818738, 1.818739, 1.81874, 1.818741, 1.818742, 1.818742, 
    1.818743, 1.818744, 1.818745, 1.818747, 1.818747, 1.818747, 1.818748, 
    1.818749, 1.818749, 1.818749, 1.818747, 1.818749, 1.818747, 1.818747, 
    1.818743, 1.818741, 1.81874, 1.81874, 1.818738, 1.818739, 1.818739, 
    1.81874, 1.818741, 1.81874, 1.818742, 1.818741, 1.818745, 1.818744, 
    1.818748, 1.818747, 1.818748, 1.818748, 1.818749, 1.818748, 1.818749, 
    1.81875, 1.818749, 1.81875, 1.818748, 1.818749, 1.81874, 1.81874, 
    1.818741, 1.81874, 1.81874, 1.818739, 1.818739, 1.81874, 1.818741, 
    1.818741, 1.818742, 1.818743, 1.818744, 1.818746, 1.818747, 1.818748, 
    1.818747, 1.818748, 1.818747, 1.818747, 1.81875, 1.818748, 1.81875, 
    1.81875, 1.818749, 1.81875, 1.81874, 1.81874, 1.818739, 1.81874, 
    1.818738, 1.818739, 1.81874, 1.818741, 1.818742, 1.818742, 1.818743, 
    1.818744, 1.818745, 1.818747, 1.818748, 1.818748, 1.818748, 1.818748, 
    1.818748, 1.818748, 1.818748, 1.818748, 1.81875, 1.81875, 1.81875, 
    1.81875, 1.81874, 1.818741, 1.81874, 1.818741, 1.818741, 1.818742, 
    1.818743, 1.818745, 1.818744, 1.818745, 1.818744, 1.818744, 1.818745, 
    1.818744, 1.818747, 1.818745, 1.818748, 1.818746, 1.818748, 1.818748, 
    1.818749, 1.818749, 1.81875, 1.818751, 1.818751, 1.818752, 1.818741, 
    1.818742, 1.818742, 1.818743, 1.818743, 1.818744, 1.818746, 1.818745, 
    1.818746, 1.818747, 1.818745, 1.818746, 1.818742, 1.818743, 1.818743, 
    1.818741, 1.818745, 1.818743, 1.818747, 1.818746, 1.818749, 1.818747, 
    1.818751, 1.818752, 1.818753, 1.818754, 1.818742, 1.818742, 1.818743, 
    1.818744, 1.818745, 1.818746, 1.818746, 1.818746, 1.818747, 1.818748, 
    1.818746, 1.818748, 1.818743, 1.818745, 1.818742, 1.818743, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818747, 1.818746, 1.818751, 1.818749, 
    1.818756, 1.818754, 1.818742, 1.818742, 1.818744, 1.818743, 1.818746, 
    1.818747, 1.818747, 1.818748, 1.818748, 1.818748, 1.818748, 1.818748, 
    1.818746, 1.818747, 1.818744, 1.818745, 1.818744, 1.818744, 1.818745, 
    1.818746, 1.818746, 1.818747, 1.818748, 1.818746, 1.818752, 1.818748, 
    1.818743, 1.818744, 1.818744, 1.818744, 1.818747, 1.818746, 1.818748, 
    1.818748, 1.818749, 1.818748, 1.818748, 1.818747, 1.818747, 1.818746, 
    1.818745, 1.818744, 1.818744, 1.818745, 1.818746, 1.818748, 1.818748, 
    1.818749, 1.818746, 1.818747, 1.818747, 1.818748, 1.818745, 1.818747, 
    1.818745, 1.818745, 1.818746, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818746, 1.818746, 1.818745, 1.818745, 1.818744, 1.818745, 
    1.818745, 1.818747, 1.818748, 1.818749, 1.818749, 1.818751, 1.81875, 
    1.818752, 1.81875, 1.818753, 1.818748, 1.81875, 1.818746, 1.818746, 
    1.818747, 1.818749, 1.818748, 1.818749, 1.818746, 1.818745, 1.818745, 
    1.818744, 1.818745, 1.818745, 1.818745, 1.818745, 1.818747, 1.818746, 
    1.818748, 1.818749, 1.818752, 1.818753, 1.818755, 1.818755, 1.818756, 
    1.818756,
  1.818756, 1.818758, 1.818758, 1.818759, 1.818758, 1.818759, 1.818757, 
    1.818758, 1.818757, 1.818756, 1.818761, 1.818759, 1.818763, 1.818762, 
    1.818766, 1.818763, 1.818766, 1.818766, 1.818767, 1.818767, 1.818769, 
    1.818768, 1.81877, 1.818769, 1.818769, 1.818768, 1.818759, 1.818761, 
    1.818759, 1.818759, 1.818759, 1.818758, 1.818758, 1.818756, 1.818756, 
    1.818757, 1.81876, 1.818759, 1.818761, 1.818761, 1.818763, 1.818762, 
    1.818765, 1.818764, 1.818767, 1.818766, 1.818767, 1.818767, 1.818767, 
    1.818766, 1.818766, 1.818765, 1.818762, 1.818763, 1.81876, 1.818758, 
    1.818757, 1.818756, 1.818756, 1.818756, 1.818757, 1.818758, 1.818759, 
    1.81876, 1.818761, 1.818762, 1.818763, 1.818765, 1.818765, 1.818766, 
    1.818766, 1.818767, 1.818767, 1.818767, 1.818766, 1.818767, 1.818765, 
    1.818765, 1.818761, 1.818759, 1.818758, 1.818758, 1.818756, 1.818757, 
    1.818757, 1.818758, 1.818758, 1.818758, 1.81876, 1.818759, 1.818763, 
    1.818762, 1.818766, 1.818765, 1.818766, 1.818766, 1.818767, 1.818766, 
    1.818768, 1.818768, 1.818768, 1.818769, 1.818766, 1.818767, 1.818758, 
    1.818758, 1.818758, 1.818757, 1.818757, 1.818756, 1.818757, 1.818757, 
    1.818758, 1.818759, 1.818759, 1.818761, 1.818762, 1.818764, 1.818765, 
    1.818766, 1.818765, 1.818766, 1.818765, 1.818765, 1.818768, 1.818766, 
    1.818769, 1.818769, 1.818767, 1.818769, 1.818758, 1.818758, 1.818757, 
    1.818758, 1.818756, 1.818757, 1.818757, 1.818759, 1.81876, 1.81876, 
    1.818761, 1.818762, 1.818763, 1.818765, 1.818766, 1.818766, 1.818766, 
    1.818766, 1.818766, 1.818767, 1.818767, 1.818766, 1.818769, 1.818768, 
    1.818769, 1.818768, 1.818758, 1.818758, 1.818758, 1.818759, 1.818758, 
    1.81876, 1.81876, 1.818763, 1.818762, 1.818763, 1.818762, 1.818762, 
    1.818763, 1.818762, 1.818765, 1.818763, 1.818766, 1.818765, 1.818767, 
    1.818766, 1.818767, 1.818767, 1.818768, 1.818769, 1.818769, 1.81877, 
    1.818759, 1.81876, 1.81876, 1.818761, 1.818761, 1.818762, 1.818764, 
    1.818763, 1.818764, 1.818765, 1.818763, 1.818764, 1.81876, 1.818761, 
    1.818761, 1.818759, 1.818763, 1.818761, 1.818765, 1.818764, 1.818767, 
    1.818766, 1.818769, 1.81877, 1.818771, 1.818773, 1.81876, 1.81876, 
    1.818761, 1.818762, 1.818763, 1.818764, 1.818764, 1.818764, 1.818765, 
    1.818766, 1.818764, 1.818766, 1.818761, 1.818763, 1.81876, 1.818761, 
    1.818762, 1.818761, 1.818763, 1.818763, 1.818765, 1.818764, 1.81877, 
    1.818767, 1.818774, 1.818772, 1.81876, 1.81876, 1.818762, 1.818761, 
    1.818764, 1.818765, 1.818765, 1.818766, 1.818766, 1.818767, 1.818766, 
    1.818767, 1.818764, 1.818765, 1.818762, 1.818763, 1.818762, 1.818762, 
    1.818763, 1.818765, 1.818765, 1.818765, 1.818766, 1.818764, 1.81877, 
    1.818766, 1.818761, 1.818762, 1.818762, 1.818762, 1.818765, 1.818764, 
    1.818767, 1.818766, 1.818767, 1.818766, 1.818766, 1.818766, 1.818765, 
    1.818764, 1.818763, 1.818762, 1.818762, 1.818763, 1.818765, 1.818766, 
    1.818766, 1.818767, 1.818764, 1.818765, 1.818765, 1.818766, 1.818763, 
    1.818766, 1.818763, 1.818763, 1.818764, 1.818765, 1.818766, 1.818766, 
    1.818766, 1.818765, 1.818764, 1.818764, 1.818763, 1.818763, 1.818762, 
    1.818763, 1.818763, 1.818765, 1.818766, 1.818767, 1.818768, 1.818769, 
    1.818768, 1.81877, 1.818768, 1.818772, 1.818766, 1.818768, 1.818764, 
    1.818764, 1.818765, 1.818767, 1.818766, 1.818767, 1.818764, 1.818763, 
    1.818763, 1.818762, 1.818763, 1.818763, 1.818763, 1.818763, 1.818765, 
    1.818764, 1.818766, 1.818767, 1.81877, 1.818772, 1.818773, 1.818774, 
    1.818774, 1.818774,
  1.818758, 1.81876, 1.818759, 1.818761, 1.81876, 1.818761, 1.818758, 
    1.81876, 1.818759, 1.818758, 1.818763, 1.818761, 1.818766, 1.818764, 
    1.818768, 1.818765, 1.818768, 1.818768, 1.818769, 1.818769, 1.818771, 
    1.81877, 1.818772, 1.818771, 1.818771, 1.81877, 1.818761, 1.818763, 
    1.818761, 1.818761, 1.818761, 1.81876, 1.818759, 1.818758, 1.818758, 
    1.818759, 1.818761, 1.818761, 1.818763, 1.818763, 1.818765, 1.818764, 
    1.818767, 1.818766, 1.818769, 1.818768, 1.818769, 1.818769, 1.818769, 
    1.818768, 1.818768, 1.818767, 1.818764, 1.818765, 1.818762, 1.81876, 
    1.818759, 1.818758, 1.818758, 1.818758, 1.818759, 1.81876, 1.818761, 
    1.818762, 1.818763, 1.818764, 1.818765, 1.818767, 1.818767, 1.818768, 
    1.818768, 1.818769, 1.818769, 1.818769, 1.818768, 1.818769, 1.818767, 
    1.818767, 1.818763, 1.818761, 1.81876, 1.81876, 1.818758, 1.818759, 
    1.818759, 1.81876, 1.81876, 1.81876, 1.818762, 1.818761, 1.818765, 
    1.818763, 1.818768, 1.818767, 1.818768, 1.818768, 1.818769, 1.818768, 
    1.81877, 1.81877, 1.81877, 1.818771, 1.818768, 1.818769, 1.81876, 
    1.81876, 1.81876, 1.818759, 1.818759, 1.818758, 1.818759, 1.818759, 
    1.81876, 1.818761, 1.818761, 1.818763, 1.818764, 1.818766, 1.818767, 
    1.818768, 1.818767, 1.818768, 1.818767, 1.818767, 1.81877, 1.818768, 
    1.818771, 1.818771, 1.818769, 1.818771, 1.81876, 1.81876, 1.818759, 
    1.818759, 1.818758, 1.818759, 1.818759, 1.818761, 1.818762, 1.818762, 
    1.818763, 1.818764, 1.818765, 1.818767, 1.818768, 1.818768, 1.818768, 
    1.818769, 1.818768, 1.818769, 1.818769, 1.818768, 1.818771, 1.81877, 
    1.818771, 1.81877, 1.81876, 1.81876, 1.81876, 1.818761, 1.81876, 
    1.818762, 1.818762, 1.818765, 1.818764, 1.818765, 1.818764, 1.818764, 
    1.818765, 1.818764, 1.818767, 1.818765, 1.818769, 1.818766, 1.818769, 
    1.818768, 1.818769, 1.818769, 1.81877, 1.818771, 1.818771, 1.818772, 
    1.818761, 1.818762, 1.818762, 1.818762, 1.818763, 1.818764, 1.818766, 
    1.818765, 1.818766, 1.818767, 1.818765, 1.818766, 1.818762, 1.818763, 
    1.818762, 1.818761, 1.818765, 1.818763, 1.818767, 1.818766, 1.818769, 
    1.818768, 1.818771, 1.818772, 1.818774, 1.818775, 1.818762, 1.818762, 
    1.818762, 1.818764, 1.818765, 1.818766, 1.818766, 1.818766, 1.818767, 
    1.818768, 1.818766, 1.818768, 1.818763, 1.818766, 1.818761, 1.818763, 
    1.818763, 1.818763, 1.818765, 1.818766, 1.818767, 1.818766, 1.818772, 
    1.818769, 1.818776, 1.818774, 1.818761, 1.818762, 1.818764, 1.818763, 
    1.818766, 1.818767, 1.818767, 1.818768, 1.818768, 1.818769, 1.818768, 
    1.818769, 1.818766, 1.818767, 1.818764, 1.818765, 1.818764, 1.818764, 
    1.818765, 1.818766, 1.818767, 1.818767, 1.818768, 1.818766, 1.818772, 
    1.818769, 1.818763, 1.818764, 1.818764, 1.818764, 1.818767, 1.818766, 
    1.818769, 1.818768, 1.818769, 1.818769, 1.818768, 1.818768, 1.818767, 
    1.818766, 1.818765, 1.818764, 1.818764, 1.818765, 1.818767, 1.818768, 
    1.818768, 1.818769, 1.818766, 1.818767, 1.818767, 1.818768, 1.818765, 
    1.818768, 1.818764, 1.818765, 1.818766, 1.818767, 1.818768, 1.818768, 
    1.818768, 1.818767, 1.818766, 1.818766, 1.818765, 1.818765, 1.818764, 
    1.818765, 1.818765, 1.818767, 1.818768, 1.818769, 1.81877, 1.818771, 
    1.81877, 1.818772, 1.81877, 1.818774, 1.818768, 1.81877, 1.818766, 
    1.818766, 1.818767, 1.818769, 1.818768, 1.818769, 1.818766, 1.818765, 
    1.818765, 1.818764, 1.818765, 1.818764, 1.818765, 1.818765, 1.818767, 
    1.818766, 1.818768, 1.818769, 1.818772, 1.818774, 1.818775, 1.818776, 
    1.818776, 1.818776,
  1.818741, 1.818742, 1.818742, 1.818743, 1.818742, 1.818743, 1.818741, 
    1.818742, 1.818741, 1.818741, 1.818745, 1.818743, 1.818748, 1.818746, 
    1.81875, 1.818748, 1.818751, 1.81875, 1.818752, 1.818751, 1.818753, 
    1.818752, 1.818755, 1.818753, 1.818753, 1.818752, 1.818744, 1.818745, 
    1.818743, 1.818744, 1.818744, 1.818742, 1.818742, 1.81874, 1.818741, 
    1.818742, 1.818744, 1.818743, 1.818745, 1.818745, 1.818747, 1.818746, 
    1.818749, 1.818748, 1.818751, 1.818751, 1.818751, 1.818751, 1.818751, 
    1.81875, 1.818751, 1.81875, 1.818746, 1.818747, 1.818744, 1.818742, 
    1.818741, 1.81874, 1.81874, 1.81874, 1.818742, 1.818743, 1.818744, 
    1.818744, 1.818745, 1.818747, 1.818748, 1.81875, 1.818749, 1.81875, 
    1.818751, 1.818751, 1.818751, 1.818752, 1.81875, 1.818751, 1.818749, 
    1.81875, 1.818745, 1.818743, 1.818743, 1.818742, 1.81874, 1.818741, 
    1.818741, 1.818742, 1.818743, 1.818742, 1.818744, 1.818743, 1.818748, 
    1.818746, 1.81875, 1.818749, 1.818751, 1.81875, 1.818751, 1.81875, 
    1.818752, 1.818752, 1.818752, 1.818753, 1.81875, 1.818751, 1.818742, 
    1.818742, 1.818743, 1.818742, 1.818741, 1.81874, 1.818741, 1.818742, 
    1.818743, 1.818743, 1.818744, 1.818745, 1.818746, 1.818748, 1.818749, 
    1.81875, 1.81875, 1.81875, 1.81875, 1.818749, 1.818752, 1.818751, 
    1.818753, 1.818753, 1.818752, 1.818753, 1.818742, 1.818742, 1.818741, 
    1.818742, 1.81874, 1.818741, 1.818742, 1.818744, 1.818744, 1.818744, 
    1.818745, 1.818746, 1.818748, 1.818749, 1.818751, 1.81875, 1.81875, 
    1.818751, 1.81875, 1.818751, 1.818751, 1.818751, 1.818753, 1.818752, 
    1.818753, 1.818752, 1.818742, 1.818743, 1.818742, 1.818743, 1.818743, 
    1.818744, 1.818745, 1.818747, 1.818746, 1.818748, 1.818746, 1.818746, 
    1.818748, 1.818746, 1.818749, 1.818747, 1.818751, 1.818749, 1.818751, 
    1.818751, 1.818751, 1.818752, 1.818752, 1.818754, 1.818753, 1.818754, 
    1.818743, 1.818744, 1.818744, 1.818745, 1.818745, 1.818746, 1.818748, 
    1.818747, 1.818749, 1.818749, 1.818747, 1.818748, 1.818745, 1.818745, 
    1.818745, 1.818743, 1.818748, 1.818745, 1.818749, 1.818748, 1.818752, 
    1.81875, 1.818753, 1.818755, 1.818756, 1.818757, 1.818744, 1.818744, 
    1.818745, 1.818746, 1.818747, 1.818748, 1.818748, 1.818749, 1.818749, 
    1.81875, 1.818749, 1.81875, 1.818745, 1.818748, 1.818744, 1.818745, 
    1.818746, 1.818745, 1.818747, 1.818748, 1.81875, 1.818749, 1.818754, 
    1.818752, 1.818758, 1.818757, 1.818744, 1.818744, 1.818747, 1.818746, 
    1.818748, 1.818749, 1.81875, 1.81875, 1.818751, 1.818751, 1.81875, 
    1.818751, 1.818748, 1.818749, 1.818746, 1.818747, 1.818747, 1.818746, 
    1.818748, 1.818749, 1.818749, 1.818749, 1.81875, 1.818748, 1.818755, 
    1.818751, 1.818745, 1.818746, 1.818746, 1.818746, 1.818749, 1.818748, 
    1.818751, 1.81875, 1.818751, 1.818751, 1.818751, 1.81875, 1.818749, 
    1.818748, 1.818747, 1.818746, 1.818746, 1.818747, 1.818749, 1.818751, 
    1.81875, 1.818751, 1.818748, 1.81875, 1.818749, 1.81875, 1.818747, 
    1.81875, 1.818747, 1.818747, 1.818748, 1.81875, 1.81875, 1.81875, 
    1.81875, 1.818749, 1.818749, 1.818748, 1.818748, 1.818747, 1.818746, 
    1.818747, 1.818748, 1.818749, 1.81875, 1.818752, 1.818752, 1.818754, 
    1.818752, 1.818755, 1.818753, 1.818756, 1.81875, 1.818753, 1.818748, 
    1.818748, 1.818749, 1.818751, 1.81875, 1.818752, 1.818749, 1.818747, 
    1.818747, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 1.818749, 
    1.818748, 1.818751, 1.818752, 1.818754, 1.818756, 1.818758, 1.818758, 
    1.818758, 1.818759,
  1.81866, 1.818661, 1.818661, 1.818662, 1.818662, 1.818662, 1.81866, 
    1.818662, 1.818661, 1.81866, 1.818664, 1.818662, 1.818667, 1.818665, 
    1.818668, 1.818666, 1.818669, 1.818668, 1.81867, 1.81867, 1.818671, 
    1.81867, 1.818673, 1.818671, 1.818671, 1.81867, 1.818663, 1.818664, 
    1.818663, 1.818663, 1.818663, 1.818662, 1.818661, 1.81866, 1.81866, 
    1.818661, 1.818663, 1.818662, 1.818664, 1.818664, 1.818666, 1.818665, 
    1.818668, 1.818667, 1.81867, 1.818669, 1.81867, 1.818669, 1.81867, 
    1.818669, 1.818669, 1.818668, 1.818665, 1.818666, 1.818663, 1.818662, 
    1.81866, 1.81866, 1.81866, 1.81866, 1.818661, 1.818662, 1.818663, 
    1.818663, 1.818664, 1.818666, 1.818666, 1.818668, 1.818668, 1.818668, 
    1.818669, 1.81867, 1.81867, 1.81867, 1.818668, 1.818669, 1.818668, 
    1.818668, 1.818664, 1.818663, 1.818662, 1.818661, 1.81866, 1.818661, 
    1.81866, 1.818661, 1.818662, 1.818662, 1.818663, 1.818663, 1.818666, 
    1.818665, 1.818669, 1.818668, 1.818669, 1.818668, 1.818669, 1.818669, 
    1.81867, 1.818671, 1.81867, 1.818671, 1.818668, 1.81867, 1.818662, 
    1.818662, 1.818662, 1.818661, 1.818661, 1.81866, 1.818661, 1.818661, 
    1.818662, 1.818663, 1.818663, 1.818664, 1.818665, 1.818667, 1.818668, 
    1.818669, 1.818668, 1.818669, 1.818668, 1.818668, 1.81867, 1.818669, 
    1.818671, 1.818671, 1.81867, 1.818671, 1.818662, 1.818661, 1.81866, 
    1.818661, 1.81866, 1.818661, 1.818661, 1.818663, 1.818663, 1.818663, 
    1.818664, 1.818665, 1.818666, 1.818668, 1.818669, 1.818669, 1.818669, 
    1.818669, 1.818668, 1.818669, 1.818669, 1.818669, 1.818671, 1.81867, 
    1.818671, 1.818671, 1.818662, 1.818662, 1.818662, 1.818662, 1.818662, 
    1.818663, 1.818664, 1.818666, 1.818665, 1.818666, 1.818665, 1.818665, 
    1.818666, 1.818665, 1.818668, 1.818666, 1.818669, 1.818667, 1.818669, 
    1.818669, 1.818669, 1.81867, 1.818671, 1.818672, 1.818671, 1.818672, 
    1.818663, 1.818663, 1.818663, 1.818664, 1.818664, 1.818665, 1.818667, 
    1.818666, 1.818667, 1.818668, 1.818666, 1.818667, 1.818664, 1.818664, 
    1.818664, 1.818663, 1.818666, 1.818664, 1.818668, 1.818667, 1.81867, 
    1.818668, 1.818671, 1.818673, 1.818674, 1.818675, 1.818664, 1.818663, 
    1.818664, 1.818665, 1.818666, 1.818667, 1.818667, 1.818667, 1.818668, 
    1.818668, 1.818667, 1.818668, 1.818664, 1.818666, 1.818663, 1.818664, 
    1.818665, 1.818664, 1.818666, 1.818667, 1.818668, 1.818667, 1.818672, 
    1.81867, 1.818676, 1.818674, 1.818663, 1.818664, 1.818665, 1.818665, 
    1.818667, 1.818668, 1.818668, 1.818669, 1.818669, 1.818669, 1.818669, 
    1.818669, 1.818667, 1.818668, 1.818665, 1.818666, 1.818666, 1.818665, 
    1.818666, 1.818667, 1.818667, 1.818668, 1.818669, 1.818667, 1.818673, 
    1.818669, 1.818664, 1.818665, 1.818665, 1.818665, 1.818668, 1.818667, 
    1.818669, 1.818669, 1.81867, 1.818669, 1.818669, 1.818668, 1.818668, 
    1.818667, 1.818666, 1.818665, 1.818665, 1.818666, 1.818668, 1.818669, 
    1.818669, 1.81867, 1.818667, 1.818668, 1.818668, 1.818669, 1.818666, 
    1.818668, 1.818666, 1.818666, 1.818667, 1.818668, 1.818668, 1.818669, 
    1.818669, 1.818668, 1.818667, 1.818667, 1.818666, 1.818666, 1.818665, 
    1.818666, 1.818666, 1.818668, 1.818669, 1.81867, 1.81867, 1.818672, 
    1.818671, 1.818673, 1.818671, 1.818674, 1.818668, 1.818671, 1.818667, 
    1.818667, 1.818668, 1.81867, 1.818669, 1.81867, 1.818667, 1.818666, 
    1.818666, 1.818665, 1.818666, 1.818666, 1.818666, 1.818666, 1.818668, 
    1.818667, 1.818669, 1.81867, 1.818672, 1.818674, 1.818675, 1.818676, 
    1.818676, 1.818676,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.592247e-09, 1.596609e-09, 1.595761e-09, 1.599278e-09, 1.597328e-09, 
    1.59963e-09, 1.593132e-09, 1.596782e-09, 1.594452e-09, 1.59264e-09, 
    1.606101e-09, 1.599435e-09, 1.613025e-09, 1.608776e-09, 1.619449e-09, 
    1.612364e-09, 1.620878e-09, 1.619246e-09, 1.62416e-09, 1.622752e-09, 
    1.629034e-09, 1.624809e-09, 1.632291e-09, 1.628026e-09, 1.628693e-09, 
    1.62467e-09, 1.600778e-09, 1.605271e-09, 1.600511e-09, 1.601152e-09, 
    1.600865e-09, 1.597368e-09, 1.595605e-09, 1.591914e-09, 1.592584e-09, 
    1.595295e-09, 1.60144e-09, 1.599355e-09, 1.604611e-09, 1.604493e-09, 
    1.610342e-09, 1.607705e-09, 1.617534e-09, 1.614741e-09, 1.622811e-09, 
    1.620782e-09, 1.622716e-09, 1.622129e-09, 1.622723e-09, 1.619747e-09, 
    1.621022e-09, 1.618403e-09, 1.608199e-09, 1.611198e-09, 1.60225e-09, 
    1.596867e-09, 1.593291e-09, 1.590754e-09, 1.591112e-09, 1.591796e-09, 
    1.595311e-09, 1.598615e-09, 1.601133e-09, 1.602817e-09, 1.604476e-09, 
    1.609494e-09, 1.612151e-09, 1.618098e-09, 1.617026e-09, 1.618843e-09, 
    1.62058e-09, 1.623494e-09, 1.623015e-09, 1.624299e-09, 1.618796e-09, 
    1.622453e-09, 1.616415e-09, 1.618066e-09, 1.604924e-09, 1.599918e-09, 
    1.597787e-09, 1.595924e-09, 1.591388e-09, 1.59452e-09, 1.593286e-09, 
    1.596224e-09, 1.59809e-09, 1.597167e-09, 1.602863e-09, 1.600649e-09, 
    1.612309e-09, 1.607287e-09, 1.620377e-09, 1.617246e-09, 1.621128e-09, 
    1.619147e-09, 1.622541e-09, 1.619487e-09, 1.624777e-09, 1.625928e-09, 
    1.625141e-09, 1.628164e-09, 1.619317e-09, 1.622715e-09, 1.597141e-09, 
    1.597291e-09, 1.597993e-09, 1.594909e-09, 1.594721e-09, 1.591895e-09, 
    1.59441e-09, 1.59548e-09, 1.598198e-09, 1.599805e-09, 1.601333e-09, 
    1.604691e-09, 1.608441e-09, 1.613683e-09, 1.617449e-09, 1.619972e-09, 
    1.618425e-09, 1.619791e-09, 1.618264e-09, 1.617549e-09, 1.625497e-09, 
    1.621034e-09, 1.62773e-09, 1.627359e-09, 1.624329e-09, 1.627401e-09, 
    1.597397e-09, 1.596531e-09, 1.593523e-09, 1.595877e-09, 1.591588e-09, 
    1.593988e-09, 1.595369e-09, 1.600694e-09, 1.601865e-09, 1.602949e-09, 
    1.605091e-09, 1.60784e-09, 1.61266e-09, 1.616854e-09, 1.620681e-09, 
    1.620401e-09, 1.620499e-09, 1.621354e-09, 1.619237e-09, 1.621702e-09, 
    1.622115e-09, 1.621034e-09, 1.62731e-09, 1.625517e-09, 1.627351e-09, 
    1.626184e-09, 1.596813e-09, 1.59827e-09, 1.597483e-09, 1.598963e-09, 
    1.59792e-09, 1.602559e-09, 1.603949e-09, 1.610455e-09, 1.607786e-09, 
    1.612034e-09, 1.608217e-09, 1.608894e-09, 1.612171e-09, 1.608424e-09, 
    1.616622e-09, 1.611064e-09, 1.621387e-09, 1.615837e-09, 1.621735e-09, 
    1.620664e-09, 1.622437e-09, 1.624024e-09, 1.626021e-09, 1.629704e-09, 
    1.628851e-09, 1.631931e-09, 1.600443e-09, 1.602333e-09, 1.602167e-09, 
    1.604145e-09, 1.605607e-09, 1.608777e-09, 1.613859e-09, 1.611948e-09, 
    1.615457e-09, 1.616161e-09, 1.610831e-09, 1.614103e-09, 1.603598e-09, 
    1.605295e-09, 1.604285e-09, 1.600592e-09, 1.612388e-09, 1.606335e-09, 
    1.617511e-09, 1.614233e-09, 1.623798e-09, 1.619041e-09, 1.628382e-09, 
    1.632372e-09, 1.636128e-09, 1.640515e-09, 1.603364e-09, 1.60208e-09, 
    1.60438e-09, 1.60756e-09, 1.610511e-09, 1.614433e-09, 1.614835e-09, 
    1.615569e-09, 1.617472e-09, 1.619072e-09, 1.615801e-09, 1.619473e-09, 
    1.605688e-09, 1.612914e-09, 1.601595e-09, 1.605003e-09, 1.607373e-09, 
    1.606334e-09, 1.61173e-09, 1.613002e-09, 1.618167e-09, 1.615497e-09, 
    1.631387e-09, 1.624359e-09, 1.643855e-09, 1.638409e-09, 1.601632e-09, 
    1.60336e-09, 1.609374e-09, 1.606513e-09, 1.614695e-09, 1.616708e-09, 
    1.618345e-09, 1.620437e-09, 1.620663e-09, 1.621902e-09, 1.619871e-09, 
    1.621822e-09, 1.614442e-09, 1.61774e-09, 1.608688e-09, 1.610891e-09, 
    1.609877e-09, 1.608765e-09, 1.612197e-09, 1.615852e-09, 1.615931e-09, 
    1.617103e-09, 1.620403e-09, 1.614728e-09, 1.632292e-09, 1.621446e-09, 
    1.605245e-09, 1.608573e-09, 1.609049e-09, 1.60776e-09, 1.616507e-09, 
    1.613338e-09, 1.621872e-09, 1.619566e-09, 1.623344e-09, 1.621466e-09, 
    1.62119e-09, 1.618779e-09, 1.617277e-09, 1.613483e-09, 1.610395e-09, 
    1.607947e-09, 1.608516e-09, 1.611206e-09, 1.616076e-09, 1.620683e-09, 
    1.619674e-09, 1.623057e-09, 1.614102e-09, 1.617857e-09, 1.616406e-09, 
    1.62019e-09, 1.611898e-09, 1.618957e-09, 1.610092e-09, 1.61087e-09, 
    1.613275e-09, 1.618111e-09, 1.619182e-09, 1.620324e-09, 1.61962e-09, 
    1.6162e-09, 1.61564e-09, 1.613217e-09, 1.612547e-09, 1.6107e-09, 
    1.609171e-09, 1.610568e-09, 1.612035e-09, 1.616202e-09, 1.619955e-09, 
    1.624046e-09, 1.625048e-09, 1.629825e-09, 1.625935e-09, 1.632352e-09, 
    1.626896e-09, 1.636341e-09, 1.619367e-09, 1.626736e-09, 1.613385e-09, 
    1.614824e-09, 1.617426e-09, 1.623393e-09, 1.620172e-09, 1.623939e-09, 
    1.615618e-09, 1.611298e-09, 1.610181e-09, 1.608095e-09, 1.610229e-09, 
    1.610055e-09, 1.612096e-09, 1.611441e-09, 1.61634e-09, 1.613709e-09, 
    1.621183e-09, 1.62391e-09, 1.631608e-09, 1.636325e-09, 1.641127e-09, 
    1.643246e-09, 1.643891e-09, 1.64416e-09 ;

 SOIL2_HR_S3 =
  1.137319e-10, 1.140435e-10, 1.139829e-10, 1.142342e-10, 1.140948e-10, 
    1.142593e-10, 1.137951e-10, 1.140558e-10, 1.138894e-10, 1.1376e-10, 
    1.147215e-10, 1.142454e-10, 1.152161e-10, 1.149125e-10, 1.15675e-10, 
    1.151688e-10, 1.15777e-10, 1.156604e-10, 1.160114e-10, 1.159109e-10, 
    1.163596e-10, 1.160578e-10, 1.165922e-10, 1.162875e-10, 1.163352e-10, 
    1.160478e-10, 1.143413e-10, 1.146622e-10, 1.143222e-10, 1.14368e-10, 
    1.143475e-10, 1.140977e-10, 1.139718e-10, 1.137081e-10, 1.13756e-10, 
    1.139496e-10, 1.143886e-10, 1.142396e-10, 1.146151e-10, 1.146066e-10, 
    1.150244e-10, 1.148361e-10, 1.155381e-10, 1.153387e-10, 1.159151e-10, 
    1.157701e-10, 1.159082e-10, 1.158664e-10, 1.159088e-10, 1.156962e-10, 
    1.157873e-10, 1.156002e-10, 1.148713e-10, 1.150856e-10, 1.144464e-10, 
    1.140619e-10, 1.138065e-10, 1.136253e-10, 1.136509e-10, 1.136997e-10, 
    1.139508e-10, 1.141868e-10, 1.143666e-10, 1.144869e-10, 1.146054e-10, 
    1.149639e-10, 1.151537e-10, 1.155784e-10, 1.155019e-10, 1.156317e-10, 
    1.157557e-10, 1.159639e-10, 1.159296e-10, 1.160213e-10, 1.156283e-10, 
    1.158895e-10, 1.154582e-10, 1.155762e-10, 1.146374e-10, 1.142798e-10, 
    1.141277e-10, 1.139946e-10, 1.136706e-10, 1.138943e-10, 1.138061e-10, 
    1.14016e-10, 1.141493e-10, 1.140834e-10, 1.144902e-10, 1.14332e-10, 
    1.151649e-10, 1.148062e-10, 1.157412e-10, 1.155176e-10, 1.157948e-10, 
    1.156534e-10, 1.158958e-10, 1.156776e-10, 1.160555e-10, 1.161377e-10, 
    1.160815e-10, 1.162975e-10, 1.156655e-10, 1.159082e-10, 1.140815e-10, 
    1.140922e-10, 1.141423e-10, 1.139221e-10, 1.139086e-10, 1.137068e-10, 
    1.138864e-10, 1.139629e-10, 1.14157e-10, 1.142718e-10, 1.143809e-10, 
    1.146208e-10, 1.148886e-10, 1.152631e-10, 1.155321e-10, 1.157123e-10, 
    1.156018e-10, 1.156994e-10, 1.155903e-10, 1.155392e-10, 1.161069e-10, 
    1.157881e-10, 1.162664e-10, 1.1624e-10, 1.160235e-10, 1.162429e-10, 
    1.140998e-10, 1.140379e-10, 1.13823e-10, 1.139912e-10, 1.136848e-10, 
    1.138563e-10, 1.139549e-10, 1.143353e-10, 1.144189e-10, 1.144964e-10, 
    1.146494e-10, 1.148457e-10, 1.1519e-10, 1.154895e-10, 1.157629e-10, 
    1.157429e-10, 1.1575e-10, 1.15811e-10, 1.156598e-10, 1.158358e-10, 
    1.158654e-10, 1.157881e-10, 1.162364e-10, 1.161084e-10, 1.162394e-10, 
    1.16156e-10, 1.14058e-10, 1.141622e-10, 1.141059e-10, 1.142117e-10, 
    1.141371e-10, 1.144685e-10, 1.145678e-10, 1.150325e-10, 1.148418e-10, 
    1.151453e-10, 1.148727e-10, 1.14921e-10, 1.151551e-10, 1.148874e-10, 
    1.15473e-10, 1.15076e-10, 1.158134e-10, 1.154169e-10, 1.158382e-10, 
    1.157617e-10, 1.158884e-10, 1.160017e-10, 1.161443e-10, 1.164074e-10, 
    1.163465e-10, 1.165665e-10, 1.143174e-10, 1.144523e-10, 1.144405e-10, 
    1.145818e-10, 1.146862e-10, 1.149126e-10, 1.152757e-10, 1.151392e-10, 
    1.153898e-10, 1.1544e-10, 1.150594e-10, 1.152931e-10, 1.145427e-10, 
    1.146639e-10, 1.145918e-10, 1.14328e-10, 1.151706e-10, 1.147382e-10, 
    1.155365e-10, 1.153024e-10, 1.159855e-10, 1.156458e-10, 1.16313e-10, 
    1.16598e-10, 1.168663e-10, 1.171796e-10, 1.14526e-10, 1.144343e-10, 
    1.145986e-10, 1.148257e-10, 1.150365e-10, 1.153167e-10, 1.153453e-10, 
    1.153978e-10, 1.155337e-10, 1.15648e-10, 1.154144e-10, 1.156766e-10, 
    1.14692e-10, 1.152081e-10, 1.143996e-10, 1.146431e-10, 1.148123e-10, 
    1.147381e-10, 1.151236e-10, 1.152144e-10, 1.155833e-10, 1.153927e-10, 
    1.165276e-10, 1.160256e-10, 1.174182e-10, 1.170292e-10, 1.144023e-10, 
    1.145257e-10, 1.149553e-10, 1.147509e-10, 1.153354e-10, 1.154792e-10, 
    1.155961e-10, 1.157455e-10, 1.157616e-10, 1.158501e-10, 1.157051e-10, 
    1.158444e-10, 1.153173e-10, 1.155529e-10, 1.149063e-10, 1.150636e-10, 
    1.149912e-10, 1.149118e-10, 1.15157e-10, 1.15418e-10, 1.154237e-10, 
    1.155073e-10, 1.157431e-10, 1.153378e-10, 1.165923e-10, 1.158176e-10, 
    1.146604e-10, 1.14898e-10, 1.14932e-10, 1.1484e-10, 1.154648e-10, 
    1.152384e-10, 1.15848e-10, 1.156833e-10, 1.159531e-10, 1.15819e-10, 
    1.157993e-10, 1.156271e-10, 1.155198e-10, 1.152488e-10, 1.150282e-10, 
    1.148533e-10, 1.14894e-10, 1.150861e-10, 1.15434e-10, 1.157631e-10, 
    1.15691e-10, 1.159326e-10, 1.15293e-10, 1.155612e-10, 1.154576e-10, 
    1.157279e-10, 1.151355e-10, 1.156398e-10, 1.150066e-10, 1.150621e-10, 
    1.152339e-10, 1.155794e-10, 1.156559e-10, 1.157374e-10, 1.156871e-10, 
    1.154428e-10, 1.154028e-10, 1.152298e-10, 1.151819e-10, 1.1505e-10, 
    1.149408e-10, 1.150406e-10, 1.151454e-10, 1.15443e-10, 1.157111e-10, 
    1.160033e-10, 1.160749e-10, 1.164161e-10, 1.161382e-10, 1.165966e-10, 
    1.162068e-10, 1.168815e-10, 1.156691e-10, 1.161954e-10, 1.152418e-10, 
    1.153445e-10, 1.155304e-10, 1.159566e-10, 1.157266e-10, 1.159957e-10, 
    1.154013e-10, 1.150927e-10, 1.150129e-10, 1.14864e-10, 1.150163e-10, 
    1.15004e-10, 1.151497e-10, 1.151029e-10, 1.154528e-10, 1.152649e-10, 
    1.157988e-10, 1.159935e-10, 1.165434e-10, 1.168804e-10, 1.172233e-10, 
    1.173747e-10, 1.174208e-10, 1.1744e-10 ;

 SOIL3C =
  5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782616, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782616, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782616, 5.782616, 
    5.782616, 5.782616 ;

 SOIL3C_TO_SOIL1C =
  3.139716e-11, 3.148315e-11, 3.146644e-11, 3.153577e-11, 3.149732e-11, 
    3.154271e-11, 3.14146e-11, 3.148655e-11, 3.144062e-11, 3.140491e-11, 
    3.167027e-11, 3.153887e-11, 3.180677e-11, 3.1723e-11, 3.193341e-11, 
    3.179373e-11, 3.196158e-11, 3.19294e-11, 3.202627e-11, 3.199852e-11, 
    3.212236e-11, 3.203908e-11, 3.218656e-11, 3.210248e-11, 3.211563e-11, 
    3.203632e-11, 3.156533e-11, 3.165391e-11, 3.156008e-11, 3.157271e-11, 
    3.156704e-11, 3.149811e-11, 3.146335e-11, 3.139059e-11, 3.14038e-11, 
    3.145725e-11, 3.157839e-11, 3.153728e-11, 3.164091e-11, 3.163856e-11, 
    3.175388e-11, 3.170189e-11, 3.189566e-11, 3.18406e-11, 3.199968e-11, 
    3.195968e-11, 3.19978e-11, 3.198624e-11, 3.199795e-11, 3.193928e-11, 
    3.196442e-11, 3.191279e-11, 3.171162e-11, 3.177075e-11, 3.159436e-11, 
    3.148823e-11, 3.141775e-11, 3.136772e-11, 3.137479e-11, 3.138827e-11, 
    3.145756e-11, 3.15227e-11, 3.157233e-11, 3.160552e-11, 3.163823e-11, 
    3.173716e-11, 3.178955e-11, 3.190678e-11, 3.188564e-11, 3.192146e-11, 
    3.19557e-11, 3.201316e-11, 3.20037e-11, 3.202901e-11, 3.192053e-11, 
    3.199262e-11, 3.187359e-11, 3.190615e-11, 3.164707e-11, 3.154838e-11, 
    3.150638e-11, 3.146965e-11, 3.138023e-11, 3.144198e-11, 3.141764e-11, 
    3.147555e-11, 3.151234e-11, 3.149415e-11, 3.160643e-11, 3.156278e-11, 
    3.179265e-11, 3.169366e-11, 3.195171e-11, 3.188998e-11, 3.19665e-11, 
    3.192746e-11, 3.199435e-11, 3.193415e-11, 3.203843e-11, 3.206113e-11, 
    3.204562e-11, 3.210522e-11, 3.193081e-11, 3.199779e-11, 3.149364e-11, 
    3.14966e-11, 3.151043e-11, 3.144964e-11, 3.144593e-11, 3.139023e-11, 
    3.14398e-11, 3.14609e-11, 3.151448e-11, 3.154616e-11, 3.157628e-11, 
    3.164248e-11, 3.17164e-11, 3.181974e-11, 3.189398e-11, 3.194373e-11, 
    3.191323e-11, 3.194016e-11, 3.191005e-11, 3.189594e-11, 3.205262e-11, 
    3.196465e-11, 3.209664e-11, 3.208935e-11, 3.202961e-11, 3.209017e-11, 
    3.149869e-11, 3.148161e-11, 3.142231e-11, 3.146872e-11, 3.138416e-11, 
    3.143149e-11, 3.14587e-11, 3.156369e-11, 3.158676e-11, 3.160814e-11, 
    3.165037e-11, 3.170455e-11, 3.179958e-11, 3.188224e-11, 3.195769e-11, 
    3.195217e-11, 3.195411e-11, 3.197096e-11, 3.192922e-11, 3.197781e-11, 
    3.198596e-11, 3.196465e-11, 3.208837e-11, 3.205303e-11, 3.208919e-11, 
    3.206618e-11, 3.148717e-11, 3.15159e-11, 3.150037e-11, 3.152956e-11, 
    3.1509e-11, 3.160044e-11, 3.162785e-11, 3.175609e-11, 3.170348e-11, 
    3.178723e-11, 3.171199e-11, 3.172532e-11, 3.178994e-11, 3.171606e-11, 
    3.187767e-11, 3.17681e-11, 3.197161e-11, 3.186221e-11, 3.197847e-11, 
    3.195737e-11, 3.199231e-11, 3.20236e-11, 3.206296e-11, 3.213556e-11, 
    3.211876e-11, 3.217947e-11, 3.155873e-11, 3.159599e-11, 3.159271e-11, 
    3.16317e-11, 3.166054e-11, 3.172302e-11, 3.182321e-11, 3.178554e-11, 
    3.18547e-11, 3.186858e-11, 3.176352e-11, 3.182802e-11, 3.162092e-11, 
    3.165438e-11, 3.163447e-11, 3.156167e-11, 3.179421e-11, 3.167488e-11, 
    3.189521e-11, 3.183059e-11, 3.201913e-11, 3.192537e-11, 3.21095e-11, 
    3.218815e-11, 3.226221e-11, 3.234868e-11, 3.161632e-11, 3.159101e-11, 
    3.163634e-11, 3.169903e-11, 3.175721e-11, 3.183453e-11, 3.184244e-11, 
    3.185692e-11, 3.189444e-11, 3.192597e-11, 3.186149e-11, 3.193387e-11, 
    3.166213e-11, 3.180457e-11, 3.158144e-11, 3.164863e-11, 3.169534e-11, 
    3.167486e-11, 3.178124e-11, 3.18063e-11, 3.190813e-11, 3.18555e-11, 
    3.216874e-11, 3.203019e-11, 3.241453e-11, 3.230717e-11, 3.158217e-11, 
    3.161624e-11, 3.17348e-11, 3.16784e-11, 3.183969e-11, 3.187938e-11, 
    3.191165e-11, 3.195287e-11, 3.195733e-11, 3.198175e-11, 3.194173e-11, 
    3.198018e-11, 3.183469e-11, 3.189972e-11, 3.172126e-11, 3.17647e-11, 
    3.174472e-11, 3.172279e-11, 3.179046e-11, 3.186251e-11, 3.186406e-11, 
    3.188716e-11, 3.195221e-11, 3.184035e-11, 3.218659e-11, 3.197278e-11, 
    3.16534e-11, 3.1719e-11, 3.172838e-11, 3.170297e-11, 3.18754e-11, 
    3.181293e-11, 3.198116e-11, 3.193571e-11, 3.201018e-11, 3.197318e-11, 
    3.196773e-11, 3.19202e-11, 3.189059e-11, 3.18158e-11, 3.175493e-11, 
    3.170666e-11, 3.171788e-11, 3.17709e-11, 3.186692e-11, 3.195773e-11, 
    3.193783e-11, 3.200452e-11, 3.1828e-11, 3.190203e-11, 3.187341e-11, 
    3.194802e-11, 3.178454e-11, 3.192371e-11, 3.174895e-11, 3.176428e-11, 
    3.181169e-11, 3.190704e-11, 3.192815e-11, 3.195066e-11, 3.193677e-11, 
    3.186935e-11, 3.185831e-11, 3.181054e-11, 3.179735e-11, 3.176094e-11, 
    3.17308e-11, 3.175834e-11, 3.178726e-11, 3.186939e-11, 3.194338e-11, 
    3.202404e-11, 3.204378e-11, 3.213795e-11, 3.206127e-11, 3.218778e-11, 
    3.20802e-11, 3.226641e-11, 3.19318e-11, 3.207706e-11, 3.181385e-11, 
    3.184222e-11, 3.189352e-11, 3.201115e-11, 3.194767e-11, 3.202192e-11, 
    3.185788e-11, 3.177273e-11, 3.17507e-11, 3.170959e-11, 3.175164e-11, 
    3.174823e-11, 3.178846e-11, 3.177553e-11, 3.187212e-11, 3.182024e-11, 
    3.196759e-11, 3.202134e-11, 3.21731e-11, 3.22661e-11, 3.236075e-11, 
    3.240252e-11, 3.241523e-11, 3.242055e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00008, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00008, 20.00009, 20.00008, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00009, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 
    20.00008, 20.00008,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256922, 0.5256923, 0.5256922, 0.5256923, 0.5256923, 0.5256923, 
    0.5256922, 0.5256923, 0.5256922, 0.5256922, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256922, 0.5256922, 0.5256922, 0.5256922, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256922, 0.5256922, 0.5256922, 0.5256922, 
    0.5256922, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256922, 0.5256922, 0.5256922, 
    0.5256922, 0.5256922, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256922, 
    0.5256922, 0.5256922, 0.5256922, 0.5256922, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256922, 0.5256922, 0.5256922, 0.5256922, 0.5256922, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  1.003089e-36, -2.569961e-21, -1.027984e-20, 2.569961e-21, -1.027984e-20, 
    -3.083953e-20, 1.541976e-20, 5.139921e-21, 5.139921e-21, 1.003089e-36, 
    -1.28498e-20, -1.28498e-20, -2.569961e-21, -2.569961e-21, -1.003089e-36, 
    -7.709882e-21, -1.027984e-20, 5.139921e-21, 0, 1.28498e-20, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -7.709882e-21, 1.28498e-20, -1.28498e-20, 2.569961e-21, -1.541976e-20, 
    1.027984e-20, 2.055969e-20, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -1.28498e-20, -1.28498e-20, -1.003089e-36, 1.541976e-20, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 1.28498e-20, 
    2.569961e-21, 1.28498e-20, 5.139921e-21, 2.055969e-20, 5.139921e-21, 
    1.003089e-36, -2.569961e-21, 2.569961e-21, 1.798972e-20, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, -5.139921e-21, 
    7.709882e-21, -7.709882e-21, 5.139921e-21, 0, 1.798972e-20, 
    -2.312965e-20, -1.027984e-20, -2.569961e-21, 2.569961e-21, 2.055969e-20, 
    -5.139921e-21, -2.055969e-20, 5.139921e-21, 1.003089e-36, 2.569961e-21, 
    1.28498e-20, 1.798972e-20, 1.28498e-20, -1.28498e-20, 5.139921e-21, 
    -1.28498e-20, 2.055969e-20, 7.709882e-21, 0, -1.027984e-20, 
    -2.312965e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -1.28498e-20, 1.28498e-20, -1.003089e-36, -1.798972e-20, -1.027984e-20, 
    5.139921e-21, -1.28498e-20, 2.055969e-20, 2.055969e-20, 0, 7.709882e-21, 
    1.798972e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, 7.709882e-21, -5.139921e-21, 0, -2.312965e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    0, 0, -1.003089e-36, 2.569961e-20, 1.28498e-20, 1.003089e-36, 
    1.003089e-36, -2.569961e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.541976e-20, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, -2.569961e-21, 1.28498e-20, 
    -1.003089e-36, 2.569961e-21, 0, -1.027984e-20, 2.569961e-21, 
    7.709882e-21, -1.003089e-36, -2.312965e-20, -7.709882e-21, 1.541976e-20, 
    1.541976e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    1.798972e-20, 7.709882e-21, 1.027984e-20, 1.28498e-20, 2.569961e-21, 
    1.28498e-20, -1.541976e-20, 1.541976e-20, 1.003089e-36, -1.003089e-36, 
    1.027984e-20, 2.055969e-20, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, 2.312965e-20, -7.709882e-21, 
    -7.709882e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, -1.003089e-36, 
    2.569961e-21, 2.569961e-21, -2.569961e-21, -1.798972e-20, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, -1.541976e-20, 2.569961e-21, 5.139921e-21, 
    1.28498e-20, 2.569961e-21, -1.003089e-36, 7.709882e-21, -7.709882e-21, 
    1.28498e-20, -2.569961e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, 1.28498e-20, -1.541976e-20, 2.569961e-21, -2.569961e-20, 
    1.027984e-20, -1.28498e-20, 1.003089e-36, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -1.541976e-20, -1.027984e-20, -5.139921e-21, 
    2.569961e-20, -2.569961e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, -1.28498e-20, -1.541976e-20, -1.28498e-20, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -1.28498e-20, 2.569961e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, -2.312965e-20, 
    1.28498e-20, 7.709882e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, 1.003089e-36, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, 1.798972e-20, 1.003089e-36, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, 1.027984e-20, 7.709882e-21, 
    1.28498e-20, -2.569961e-21, 1.28498e-20, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-20, -2.312965e-20, -1.541976e-20, 1.541976e-20, 
    1.541976e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 
    -7.709882e-21, 1.003089e-36, -2.055969e-20, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, -2.055969e-20, 
    1.027984e-20, 7.709882e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -1.798972e-20, -1.541976e-20, 1.28498e-20, -2.569961e-21, 
    2.312965e-20, -1.003089e-36, 7.709882e-21, -5.139921e-21, -1.798972e-20, 
    -1.28498e-20, 7.709882e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, -5.139921e-21, 1.003089e-36, 
    2.569961e-21, 1.798972e-20, 2.569961e-21, -1.541976e-20, -2.569961e-21, 
    -2.569961e-21, 0, 7.709882e-21, 5.139921e-21, 7.709882e-21, 
    -1.541976e-20, 1.027984e-20, 1.28498e-20, 2.569961e-21, 0, -2.569961e-21, 
    -1.28498e-20, -7.709882e-21, -1.541976e-20, 7.709882e-21, 2.569961e-21, 
    1.027984e-20,
  0, -1.027984e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, -7.709882e-21, 
    -1.28498e-20, 2.569961e-21, 0, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 0, -7.709882e-21, 1.027984e-20, -1.027984e-20, 
    7.709882e-21, -1.003089e-36, -1.28498e-20, 1.003089e-36, -2.055969e-20, 
    1.28498e-20, -7.709882e-21, 2.569961e-21, 0, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 7.709882e-21, 1.003089e-36, 0, 
    5.139921e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, 0, 2.569961e-21, -2.569961e-21, 
    1.541976e-20, -1.027984e-20, -1.28498e-20, 2.569961e-21, -1.541976e-20, 
    -2.569961e-21, 5.139921e-21, -7.709882e-21, 1.027984e-20, -1.003089e-36, 
    -1.541976e-20, -2.569961e-21, 0, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, 1.027984e-20, 1.027984e-20, -7.709882e-21, -1.027984e-20, 
    2.569961e-21, 0, -1.027984e-20, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -1.027984e-20, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, 5.139921e-21, 
    0, 2.569961e-21, 0, -1.28498e-20, 1.027984e-20, 0, -7.709882e-21, 
    1.027984e-20, -1.003089e-36, 0, -2.569961e-21, -2.569961e-21, 
    -1.28498e-20, -7.709882e-21, 0, 2.569961e-21, 1.798972e-20, 7.709882e-21, 
    1.027984e-20, -1.003089e-36, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -1.28498e-20, -1.027984e-20, 2.569961e-21, 2.569961e-21, 7.709882e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 0, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, -1.798972e-20, 5.139921e-21, 
    -2.569961e-21, 0, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, -1.027984e-20, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 1.003089e-36, 1.798972e-20, 
    2.569961e-21, -1.027984e-20, -5.139921e-21, -1.28498e-20, 2.569961e-21, 
    -2.569961e-21, 0, 0, -7.709882e-21, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    0, 5.139921e-21, -1.28498e-20, -2.569961e-21, -7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, 2.569961e-21, 0, 2.569961e-21, 1.28498e-20, 
    1.027984e-20, 1.28498e-20, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    2.569961e-21, -2.312965e-20, 2.569961e-21, 1.28498e-20, 0, -2.569961e-21, 
    0, 2.569961e-21, 7.709882e-21, -2.569961e-21, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, -1.027984e-20, 
    2.569961e-21, 2.569961e-21, -1.003089e-36, 0, -7.709882e-21, 1.28498e-20, 
    -7.709882e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, 1.003089e-36, 1.027984e-20, -7.709882e-21, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, 1.027984e-20, -1.28498e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 0, 
    -7.709882e-21, 7.709882e-21, 0, 1.027984e-20, 1.541976e-20, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 0, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, -1.28498e-20, -1.541976e-20, 
    2.569961e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    1.28498e-20, 2.569961e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, 1.28498e-20, 7.709882e-21, -1.027984e-20, 
    1.003089e-36, -5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 0, 
    0, 2.569961e-21, -7.709882e-21, -7.709882e-21, 1.541976e-20, 
    -1.027984e-20, 1.28498e-20, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -5.139921e-21, 0, 7.709882e-21, -5.139921e-21, 
    1.003089e-36, 1.003089e-36, 2.569961e-21, -7.709882e-21, 7.709882e-21, 
    7.709882e-21, 2.569961e-21, 1.28498e-20, 7.709882e-21, -1.027984e-20, 
    2.569961e-21, -1.798972e-20, -5.139921e-21, -5.139921e-21, 7.709882e-21, 
    7.709882e-21, -1.027984e-20, 0, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, 0, -1.027984e-20, 1.798972e-20, -7.709882e-21, 
    5.139921e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 
    -7.709882e-21, 0, -2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -5.139921e-21, -1.28498e-20, 5.139921e-21, 2.569961e-21, -1.28498e-20, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 1.003089e-36, 
    2.569961e-21, -1.003089e-36, 0, 0,
  -2.569961e-21, 1.798972e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -1.541976e-20, -7.709882e-21, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    1.027984e-20, 1.027984e-20, -2.569961e-21, -1.003089e-36, 0, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, -2.569961e-21, 1.28498e-20, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 1.003089e-36, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    -2.569961e-21, 2.569961e-21, -1.28498e-20, -1.28498e-20, 5.139921e-21, 
    2.569961e-20, -1.003089e-36, 0, 1.027984e-20, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 0, -7.709882e-21, 2.569961e-21, 
    -1.541976e-20, 5.139921e-21, -7.709882e-21, 1.541976e-20, 1.003089e-36, 
    1.28498e-20, 1.027984e-20, 5.139921e-21, -7.709882e-21, 1.027984e-20, 
    2.569961e-21, 1.28498e-20, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -7.709882e-21, 0, 7.709882e-21, 0, -1.027984e-20, 2.569961e-21, 0, 
    7.709882e-21, -1.28498e-20, 7.709882e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -2.055969e-20, 1.027984e-20, 2.569961e-21, 7.709882e-21, 
    1.027984e-20, 0, -5.139921e-21, -1.541976e-20, -1.28498e-20, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, 1.541976e-20, 0, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -1.027984e-20, -7.709882e-21, 1.28498e-20, 5.139921e-21, 5.139921e-21, 
    -1.28498e-20, -7.709882e-21, 1.003089e-36, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 0, 0, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, 1.027984e-20, 0, -2.569961e-21, 1.003089e-36, 
    -1.027984e-20, -7.709882e-21, 1.003089e-36, 0, 3.083953e-20, 
    1.027984e-20, 1.28498e-20, -2.569961e-21, -1.798972e-20, 1.003089e-36, 
    -1.003089e-36, 1.003089e-36, 2.569961e-21, -1.541976e-20, 1.28498e-20, 
    7.709882e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    5.139921e-21, -1.541976e-20, -1.027984e-20, 0, -2.569961e-21, 
    1.28498e-20, 1.027984e-20, -5.139921e-21, 0, -5.139921e-21, 1.003089e-36, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, -7.709882e-21, 0, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -1.28498e-20, 1.28498e-20, -1.003089e-36, 1.541976e-20, 
    -1.28498e-20, 7.709882e-21, 1.28498e-20, 1.28498e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, 0, 5.139921e-21, 2.569961e-21, 
    -1.28498e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.28498e-20, -5.139921e-21, 0, 1.798972e-20, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, 1.541976e-20, 
    -5.139921e-21, 1.003089e-36, 1.003089e-36, 1.541976e-20, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, -7.709882e-21, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 0, 
    1.28498e-20, 5.139921e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, 0, 0, -1.541976e-20, -1.541976e-20, -7.709882e-21, 
    -1.28498e-20, 1.027984e-20, 0, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -2.055969e-20, 1.027984e-20, -7.709882e-21, -5.139921e-21, 
    7.709882e-21, -1.003089e-36, -1.541976e-20, -1.027984e-20, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, -1.003089e-36, 
    0, -2.569961e-21, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, -1.541976e-20, 1.798972e-20, 0, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, 0, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, -1.027984e-20, -7.709882e-21, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 0, -7.709882e-21, 
    -1.003089e-36, -7.709882e-21, 1.027984e-20, -2.569961e-21, 1.027984e-20, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -1.541976e-20, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, -2.569961e-21, 0, 
    1.541976e-20, 7.709882e-21, 0, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -1.003089e-36, -2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21,
  -1.027984e-20, -2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-20, -1.027984e-20, -1.003089e-36, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    1.28498e-20, 0, 1.541976e-20, -1.003089e-36, 1.003089e-36, -7.709882e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 1.28498e-20, 1.027984e-20, -1.541976e-20, 
    -7.709882e-21, -5.139921e-21, 2.569961e-20, 5.139921e-21, 5.139921e-21, 
    0, 5.139921e-21, -2.569961e-21, 2.569961e-20, 2.055969e-20, 
    -2.569961e-21, -1.28498e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, 7.709882e-21, -1.027984e-20, -7.709882e-21, -1.798972e-20, 
    -1.003089e-36, 2.569961e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 7.709882e-21, -1.28498e-20, -3.083953e-20, 
    -1.541976e-20, 0, -7.709882e-21, 5.139921e-21, 1.027984e-20, 
    2.312965e-20, 2.569961e-21, -2.569961e-21, -7.709882e-21, -7.709882e-21, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, -1.798972e-20, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, -1.027984e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, -1.798972e-20, 7.709882e-21, 
    -1.003089e-36, 1.027984e-20, -2.569961e-21, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, -7.709882e-21, -1.027984e-20, 
    1.003089e-36, 1.027984e-20, -2.569961e-21, 2.569961e-21, 1.003089e-36, 
    -2.569961e-21, -1.28498e-20, -5.139921e-21, 7.709882e-21, -1.28498e-20, 
    7.709882e-21, 1.28498e-20, 1.027984e-20, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 0, 1.28498e-20, -5.139921e-21, -2.569961e-20, 0, 
    1.541976e-20, -1.027984e-20, -2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -1.003089e-36, 2.569961e-21, 0, 
    -5.139921e-21, 5.139921e-21, 1.28498e-20, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -1.28498e-20, -1.798972e-20, 
    -7.709882e-21, -1.027984e-20, 0, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, -1.28498e-20, 1.28498e-20, 2.569961e-21, 1.027984e-20, 
    1.027984e-20, -7.709882e-21, -1.027984e-20, 2.569961e-21, 1.027984e-20, 
    0, -7.709882e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -1.28498e-20, 7.709882e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, 
    1.28498e-20, -1.003089e-36, -1.541976e-20, -1.027984e-20, 0, 
    -1.28498e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, 0, 0, -1.027984e-20, 1.027984e-20, 
    7.709882e-21, -1.003089e-36, -1.28498e-20, 1.027984e-20, 1.027984e-20, 
    -1.003089e-36, 5.139921e-21, 2.569961e-20, -7.709882e-21, 1.003089e-36, 
    -1.28498e-20, -5.139921e-21, -7.709882e-21, 0, 1.28498e-20, -1.28498e-20, 
    7.709882e-21, -2.569961e-21, 1.28498e-20, 1.798972e-20, -1.027984e-20, 
    5.139921e-21, -2.569961e-21, 1.541976e-20, 7.709882e-21, 1.28498e-20, 
    -7.709882e-21, 5.139921e-21, -7.709882e-21, -2.055969e-20, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, 2.569961e-21, 1.28498e-20, 7.709882e-21, 
    -1.027984e-20, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, 5.139921e-21, -2.569961e-20, 
    -1.541976e-20, -1.027984e-20, 0, -7.709882e-21, -2.569961e-21, 
    1.28498e-20, 2.569961e-21, -2.569961e-21, 1.541976e-20, 7.709882e-21, 
    -1.027984e-20, 2.055969e-20, -5.139921e-21, 5.139921e-21, 2.055969e-20, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, -1.798972e-20, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 
    1.003089e-36, -2.569961e-21, -1.798972e-20, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 1.798972e-20, 2.569961e-21, -1.003089e-36, 1.28498e-20, 
    -2.569961e-21, 5.139921e-21, -1.003089e-36, 2.569961e-21, -1.28498e-20, 
    -2.312965e-20, -1.798972e-20, -1.28498e-20, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.541976e-20, -7.709882e-21, -7.709882e-21, 
    -5.139921e-21, -1.003089e-36, -7.709882e-21, 1.003089e-36, -1.027984e-20, 
    2.569961e-21, 5.139921e-21, 1.28498e-20, -5.139921e-21, 1.798972e-20, 
    1.003089e-36, 5.139921e-21, 2.569961e-21, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 1.28498e-20, -7.709882e-21, 
    7.709882e-21, 2.569961e-21, 2.312965e-20, 1.798972e-20, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, 2.055969e-20, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, -1.541976e-20, -2.569961e-21, 1.798972e-20, 1.027984e-20, 
    2.569961e-21, 2.569961e-20, -1.798972e-20, -1.027984e-20, 7.709882e-21, 
    7.709882e-21, 7.709882e-21, -7.709882e-21, 1.027984e-20, -1.28498e-20, 
    -1.003089e-36, -3.340949e-20, -5.139921e-21, -1.027984e-20, 
    -1.798972e-20, -5.139921e-21,
  1.003089e-36, -2.569961e-21, -2.569961e-21, -1.798972e-20, 5.139921e-21, 
    2.569961e-21, 1.798972e-20, 7.709882e-21, 1.541976e-20, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, -5.139921e-21, 1.798972e-20, -1.541976e-20, 
    1.003089e-36, -1.027984e-20, -7.709882e-21, 1.027984e-20, 2.826957e-20, 
    1.003089e-36, -1.28498e-20, -2.569961e-21, 2.055969e-20, -1.798972e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -1.027984e-20, 2.055969e-20, -2.055969e-20, 2.569961e-21, 
    1.027984e-20, 0, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, 1.003089e-36, -1.28498e-20, 
    -5.139921e-21, 2.569961e-21, 0, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 0, 2.055969e-20, -2.569961e-21, 0, -1.003089e-36, 
    -5.139921e-21, 2.569961e-20, 0, 1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 5.139921e-21, -7.709882e-21, 
    2.055969e-20, 7.709882e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 1.003089e-36, 7.709882e-21, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 1.28498e-20, 0, -5.139921e-21, -7.709882e-21, 
    -1.28498e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, 1.003089e-36, 
    -5.015443e-37, 5.139921e-21, -2.569961e-21, 0, -1.28498e-20, 
    -1.798972e-20, -1.027984e-20, 2.569961e-21, -5.139921e-21, 1.541976e-20, 
    1.027984e-20, 2.569961e-21, 1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -1.027984e-20, -2.055969e-20, -7.709882e-21, 1.027984e-20, -5.139921e-21, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, -1.28498e-20, 
    7.709882e-21, -1.003089e-36, -7.709882e-21, 1.541976e-20, -1.798972e-20, 
    1.541976e-20, -1.027984e-20, 1.28498e-20, -2.569961e-21, 1.541976e-20, 
    1.541976e-20, -7.709882e-21, -2.569961e-21, -2.312965e-20, -1.027984e-20, 
    2.569961e-21, 0, 7.709882e-21, 3.009266e-36, 3.597945e-20, 7.709882e-21, 
    -1.027984e-20, 1.798972e-20, 1.28498e-20, 1.28498e-20, 1.027984e-20, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, 7.709882e-21, -1.798972e-20, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-21, -1.798972e-20, 
    -2.055969e-20, 2.569961e-21, 7.709882e-21, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, 0, -5.139921e-21, -1.003089e-36, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -1.027984e-20, 1.003089e-36, -1.541976e-20, 
    1.28498e-20, 1.003089e-36, 0, 7.709882e-21, -2.569961e-21, 1.003089e-36, 
    -1.003089e-36, -1.003089e-36, -1.28498e-20, 5.139921e-21, 1.28498e-20, 
    5.139921e-21, 5.139921e-21, 1.798972e-20, -2.569961e-21, 1.003089e-36, 
    -5.139921e-21, -1.28498e-20, 1.28498e-20, -1.003089e-36, 1.027984e-20, 
    1.798972e-20, -7.709882e-21, -1.541976e-20, 1.28498e-20, -2.569961e-21, 
    5.139921e-21, 1.003089e-36, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    1.28498e-20, 7.709882e-21, -1.541976e-20, 0, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, -1.28498e-20, 1.28498e-20, 7.709882e-21, 7.709882e-21, 
    -1.027984e-20, 1.027984e-20, 2.569961e-21, 1.28498e-20, 7.709882e-21, 
    -5.139921e-21, 1.798972e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    1.027984e-20, -1.28498e-20, 2.569961e-21, 1.28498e-20, 1.003089e-36, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, -1.027984e-20, 
    -7.709882e-21, -7.709882e-21, -1.027984e-20, -7.709882e-21, 7.709882e-21, 
    2.569961e-21, 2.055969e-20, 1.027984e-20, 0, -1.798972e-20, 1.027984e-20, 
    -1.541976e-20, 5.139921e-21, 7.709882e-21, -1.027984e-20, -1.541976e-20, 
    -7.709882e-21, 0, 1.541976e-20, 1.28498e-20, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, -1.003089e-36, 2.569961e-21, 
    -2.312965e-20, 7.709882e-21, -1.798972e-20, -2.569961e-21, -7.709882e-21, 
    -2.312965e-20, 1.003089e-36, 5.139921e-21, -1.28498e-20, -5.139921e-21, 
    -1.027984e-20, -1.28498e-20, 2.569961e-21, 1.28498e-20, -2.569961e-21, 
    1.798972e-20, 2.569961e-21, -1.003089e-36, 5.139921e-21, -7.709882e-21, 
    2.569961e-20, 1.003089e-36, 1.28498e-20, -2.569961e-21, 1.027984e-20, 
    -1.027984e-20, -2.569961e-21, -1.541976e-20, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, -1.28498e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 
    -1.798972e-20, 5.139921e-21, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    1.28498e-20, 1.027984e-20, -1.798972e-20, -1.541976e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-20, 2.055969e-20, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, -1.28498e-20, 1.28498e-20, 
    -1.027984e-20, 7.709882e-21, -2.569961e-21, -1.798972e-20, 2.569961e-21, 
    2.569961e-21, -1.798972e-20, 2.569961e-21, -7.709882e-21, 2.569961e-20, 
    5.139921e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, 1.28498e-20, 
    -1.28498e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 1.798972e-20, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 1.541976e-20,
  6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.25807e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.25807e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  6.34286e-12, 6.360231e-12, 6.356856e-12, 6.370863e-12, 6.363094e-12, 
    6.372265e-12, 6.346383e-12, 6.36092e-12, 6.351641e-12, 6.344425e-12, 
    6.398034e-12, 6.371488e-12, 6.42561e-12, 6.408686e-12, 6.451195e-12, 
    6.422975e-12, 6.456884e-12, 6.450384e-12, 6.469953e-12, 6.464348e-12, 
    6.489366e-12, 6.47254e-12, 6.502335e-12, 6.48535e-12, 6.488006e-12, 
    6.471985e-12, 6.376834e-12, 6.394729e-12, 6.375773e-12, 6.378325e-12, 
    6.37718e-12, 6.363254e-12, 6.356232e-12, 6.341534e-12, 6.344203e-12, 
    6.354999e-12, 6.379473e-12, 6.371168e-12, 6.392102e-12, 6.391629e-12, 
    6.414925e-12, 6.404423e-12, 6.443567e-12, 6.432444e-12, 6.464582e-12, 
    6.456501e-12, 6.464202e-12, 6.461867e-12, 6.464232e-12, 6.45238e-12, 
    6.457458e-12, 6.447029e-12, 6.406389e-12, 6.418334e-12, 6.382699e-12, 
    6.361259e-12, 6.34702e-12, 6.336913e-12, 6.338342e-12, 6.341065e-12, 
    6.355063e-12, 6.368222e-12, 6.378249e-12, 6.384954e-12, 6.391561e-12, 
    6.411548e-12, 6.422131e-12, 6.445814e-12, 6.441543e-12, 6.44878e-12, 
    6.455697e-12, 6.467304e-12, 6.465395e-12, 6.470507e-12, 6.448591e-12, 
    6.463156e-12, 6.43911e-12, 6.445687e-12, 6.393348e-12, 6.373409e-12, 
    6.364925e-12, 6.357504e-12, 6.339441e-12, 6.351915e-12, 6.346998e-12, 
    6.358697e-12, 6.36613e-12, 6.362454e-12, 6.385138e-12, 6.37632e-12, 
    6.422757e-12, 6.402759e-12, 6.45489e-12, 6.44242e-12, 6.457879e-12, 
    6.449992e-12, 6.463505e-12, 6.451343e-12, 6.472411e-12, 6.476996e-12, 
    6.473863e-12, 6.485903e-12, 6.450669e-12, 6.464201e-12, 6.362351e-12, 
    6.362951e-12, 6.365743e-12, 6.353464e-12, 6.352713e-12, 6.34146e-12, 
    6.351474e-12, 6.355737e-12, 6.366561e-12, 6.372962e-12, 6.379046e-12, 
    6.39242e-12, 6.407353e-12, 6.428231e-12, 6.443228e-12, 6.453278e-12, 
    6.447117e-12, 6.452556e-12, 6.446475e-12, 6.443625e-12, 6.475277e-12, 
    6.457505e-12, 6.484171e-12, 6.482696e-12, 6.470629e-12, 6.482862e-12, 
    6.363371e-12, 6.359922e-12, 6.347941e-12, 6.357317e-12, 6.340234e-12, 
    6.349796e-12, 6.355293e-12, 6.376502e-12, 6.381163e-12, 6.385482e-12, 
    6.394014e-12, 6.404959e-12, 6.424157e-12, 6.440857e-12, 6.4561e-12, 
    6.454983e-12, 6.455376e-12, 6.45878e-12, 6.450347e-12, 6.460164e-12, 
    6.461811e-12, 6.457504e-12, 6.482499e-12, 6.475359e-12, 6.482665e-12, 
    6.478016e-12, 6.361044e-12, 6.366848e-12, 6.363712e-12, 6.369609e-12, 
    6.365454e-12, 6.383927e-12, 6.389465e-12, 6.415373e-12, 6.404744e-12, 
    6.421662e-12, 6.406463e-12, 6.409156e-12, 6.42221e-12, 6.407285e-12, 
    6.439934e-12, 6.417798e-12, 6.458912e-12, 6.436809e-12, 6.460297e-12, 
    6.456034e-12, 6.463093e-12, 6.469413e-12, 6.477366e-12, 6.492033e-12, 
    6.488637e-12, 6.500904e-12, 6.375501e-12, 6.383027e-12, 6.382366e-12, 
    6.390243e-12, 6.396067e-12, 6.408691e-12, 6.428932e-12, 6.421322e-12, 
    6.435293e-12, 6.438097e-12, 6.416872e-12, 6.429903e-12, 6.388065e-12, 
    6.394825e-12, 6.390802e-12, 6.376094e-12, 6.423073e-12, 6.398967e-12, 
    6.443476e-12, 6.430422e-12, 6.468511e-12, 6.44957e-12, 6.486768e-12, 
    6.502658e-12, 6.517618e-12, 6.535087e-12, 6.387136e-12, 6.382023e-12, 
    6.391181e-12, 6.403845e-12, 6.415599e-12, 6.431218e-12, 6.432817e-12, 
    6.435742e-12, 6.44332e-12, 6.449691e-12, 6.436665e-12, 6.451287e-12, 
    6.396389e-12, 6.425166e-12, 6.380088e-12, 6.393663e-12, 6.403099e-12, 
    6.398962e-12, 6.420453e-12, 6.425516e-12, 6.446087e-12, 6.435455e-12, 
    6.498735e-12, 6.470746e-12, 6.54839e-12, 6.5267e-12, 6.380236e-12, 
    6.38712e-12, 6.41107e-12, 6.399676e-12, 6.432261e-12, 6.440279e-12, 
    6.446797e-12, 6.455126e-12, 6.456026e-12, 6.460961e-12, 6.452875e-12, 
    6.460642e-12, 6.431251e-12, 6.444387e-12, 6.408335e-12, 6.417111e-12, 
    6.413074e-12, 6.408646e-12, 6.422314e-12, 6.43687e-12, 6.437184e-12, 
    6.44185e-12, 6.454991e-12, 6.432394e-12, 6.502341e-12, 6.459148e-12, 
    6.394626e-12, 6.407878e-12, 6.409774e-12, 6.40464e-12, 6.439475e-12, 
    6.426855e-12, 6.460841e-12, 6.451658e-12, 6.466704e-12, 6.459228e-12, 
    6.458127e-12, 6.448524e-12, 6.442544e-12, 6.427433e-12, 6.415136e-12, 
    6.405385e-12, 6.407653e-12, 6.418364e-12, 6.437761e-12, 6.456106e-12, 
    6.452088e-12, 6.46556e-12, 6.4299e-12, 6.444854e-12, 6.439074e-12, 
    6.454145e-12, 6.421119e-12, 6.449235e-12, 6.413929e-12, 6.417026e-12, 
    6.426605e-12, 6.445866e-12, 6.450131e-12, 6.454679e-12, 6.451873e-12, 
    6.438254e-12, 6.436023e-12, 6.426372e-12, 6.423706e-12, 6.416352e-12, 
    6.410262e-12, 6.415826e-12, 6.421668e-12, 6.43826e-12, 6.453209e-12, 
    6.469502e-12, 6.473491e-12, 6.492515e-12, 6.477025e-12, 6.502581e-12, 
    6.480849e-12, 6.518467e-12, 6.450868e-12, 6.480214e-12, 6.427042e-12, 
    6.432773e-12, 6.443135e-12, 6.4669e-12, 6.454074e-12, 6.469075e-12, 
    6.435936e-12, 6.418732e-12, 6.414284e-12, 6.405978e-12, 6.414474e-12, 
    6.413783e-12, 6.421912e-12, 6.4193e-12, 6.438811e-12, 6.428331e-12, 
    6.458099e-12, 6.468958e-12, 6.499617e-12, 6.518403e-12, 6.537525e-12, 
    6.545964e-12, 6.548532e-12, 6.549606e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 1.81819, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819,
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 
    1.818189, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 
    1.818189, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.83743e-11, 3.84794e-11, 3.845898e-11, 3.854372e-11, 3.849672e-11, 
    3.85522e-11, 3.839562e-11, 3.848356e-11, 3.842743e-11, 3.838378e-11, 
    3.870811e-11, 3.854751e-11, 3.887494e-11, 3.877255e-11, 3.902973e-11, 
    3.8859e-11, 3.906415e-11, 3.902483e-11, 3.914322e-11, 3.910931e-11, 
    3.926066e-11, 3.915887e-11, 3.933913e-11, 3.923637e-11, 3.925243e-11, 
    3.915551e-11, 3.857985e-11, 3.868811e-11, 3.857343e-11, 3.858887e-11, 
    3.858194e-11, 3.849768e-11, 3.84552e-11, 3.836628e-11, 3.838243e-11, 
    3.844775e-11, 3.859581e-11, 3.854557e-11, 3.867221e-11, 3.866936e-11, 
    3.88103e-11, 3.874676e-11, 3.898358e-11, 3.891629e-11, 3.911072e-11, 
    3.906183e-11, 3.910842e-11, 3.90943e-11, 3.910861e-11, 3.90369e-11, 
    3.906762e-11, 3.900453e-11, 3.875865e-11, 3.883092e-11, 3.861533e-11, 
    3.848561e-11, 3.839947e-11, 3.833832e-11, 3.834697e-11, 3.836344e-11, 
    3.844813e-11, 3.852775e-11, 3.858841e-11, 3.862898e-11, 3.866895e-11, 
    3.878986e-11, 3.885389e-11, 3.899717e-11, 3.897134e-11, 3.901512e-11, 
    3.905697e-11, 3.912719e-11, 3.911564e-11, 3.914657e-11, 3.901398e-11, 
    3.91021e-11, 3.895661e-11, 3.899641e-11, 3.867975e-11, 3.855913e-11, 
    3.850779e-11, 3.84629e-11, 3.835362e-11, 3.842908e-11, 3.839934e-11, 
    3.847012e-11, 3.851509e-11, 3.849285e-11, 3.863008e-11, 3.857674e-11, 
    3.885768e-11, 3.873669e-11, 3.905208e-11, 3.897664e-11, 3.907017e-11, 
    3.902245e-11, 3.910421e-11, 3.903063e-11, 3.915809e-11, 3.918583e-11, 
    3.916687e-11, 3.923971e-11, 3.902655e-11, 3.910841e-11, 3.849222e-11, 
    3.849585e-11, 3.851275e-11, 3.843846e-11, 3.843391e-11, 3.836583e-11, 
    3.842641e-11, 3.845221e-11, 3.85177e-11, 3.855642e-11, 3.859323e-11, 
    3.867414e-11, 3.876449e-11, 3.88908e-11, 3.898153e-11, 3.904233e-11, 
    3.900506e-11, 3.903797e-11, 3.900117e-11, 3.898393e-11, 3.917543e-11, 
    3.906791e-11, 3.922923e-11, 3.922031e-11, 3.91473e-11, 3.922132e-11, 
    3.84984e-11, 3.847753e-11, 3.840504e-11, 3.846177e-11, 3.835842e-11, 
    3.841627e-11, 3.844952e-11, 3.857784e-11, 3.860604e-11, 3.863217e-11, 
    3.868378e-11, 3.875001e-11, 3.886615e-11, 3.896718e-11, 3.90594e-11, 
    3.905265e-11, 3.905503e-11, 3.907562e-11, 3.90246e-11, 3.908399e-11, 
    3.909395e-11, 3.90679e-11, 3.921911e-11, 3.917592e-11, 3.922012e-11, 
    3.9192e-11, 3.848431e-11, 3.851943e-11, 3.850045e-11, 3.853614e-11, 
    3.851099e-11, 3.862276e-11, 3.865626e-11, 3.8813e-11, 3.87487e-11, 
    3.885106e-11, 3.87591e-11, 3.87754e-11, 3.885437e-11, 3.876408e-11, 
    3.89616e-11, 3.882768e-11, 3.907642e-11, 3.89427e-11, 3.908479e-11, 
    3.9059e-11, 3.910171e-11, 3.913995e-11, 3.918806e-11, 3.92768e-11, 
    3.925626e-11, 3.933047e-11, 3.857178e-11, 3.861731e-11, 3.861332e-11, 
    3.866097e-11, 3.869621e-11, 3.877258e-11, 3.889504e-11, 3.8849e-11, 
    3.893353e-11, 3.895049e-11, 3.882207e-11, 3.890091e-11, 3.86478e-11, 
    3.868869e-11, 3.866435e-11, 3.857537e-11, 3.885959e-11, 3.871375e-11, 
    3.898303e-11, 3.890405e-11, 3.913449e-11, 3.90199e-11, 3.924494e-11, 
    3.934108e-11, 3.943159e-11, 3.953728e-11, 3.864218e-11, 3.861124e-11, 
    3.866664e-11, 3.874326e-11, 3.881437e-11, 3.890887e-11, 3.891854e-11, 
    3.893624e-11, 3.898209e-11, 3.902063e-11, 3.894183e-11, 3.903029e-11, 
    3.869816e-11, 3.887225e-11, 3.859953e-11, 3.868166e-11, 3.873875e-11, 
    3.871372e-11, 3.884374e-11, 3.887437e-11, 3.899883e-11, 3.89345e-11, 
    3.931734e-11, 3.914801e-11, 3.961776e-11, 3.948654e-11, 3.860042e-11, 
    3.864208e-11, 3.878698e-11, 3.871804e-11, 3.891518e-11, 3.896369e-11, 
    3.900312e-11, 3.905351e-11, 3.905896e-11, 3.908881e-11, 3.903989e-11, 
    3.908688e-11, 3.890907e-11, 3.898854e-11, 3.877043e-11, 3.882352e-11, 
    3.87991e-11, 3.87723e-11, 3.8855e-11, 3.894306e-11, 3.894496e-11, 
    3.897319e-11, 3.90527e-11, 3.891598e-11, 3.933916e-11, 3.907785e-11, 
    3.868748e-11, 3.876766e-11, 3.877913e-11, 3.874807e-11, 3.895882e-11, 
    3.888247e-11, 3.908809e-11, 3.903253e-11, 3.912356e-11, 3.907833e-11, 
    3.907167e-11, 3.901357e-11, 3.897739e-11, 3.888597e-11, 3.881158e-11, 
    3.875258e-11, 3.87663e-11, 3.88311e-11, 3.894845e-11, 3.905944e-11, 
    3.903513e-11, 3.911664e-11, 3.890089e-11, 3.899137e-11, 3.895639e-11, 
    3.904758e-11, 3.884777e-11, 3.901787e-11, 3.880427e-11, 3.882301e-11, 
    3.888096e-11, 3.899749e-11, 3.902329e-11, 3.905081e-11, 3.903383e-11, 
    3.895144e-11, 3.893794e-11, 3.887955e-11, 3.886342e-11, 3.881893e-11, 
    3.878208e-11, 3.881575e-11, 3.885109e-11, 3.895147e-11, 3.904191e-11, 
    3.914049e-11, 3.916462e-11, 3.927971e-11, 3.9186e-11, 3.934061e-11, 
    3.920914e-11, 3.943672e-11, 3.902775e-11, 3.92053e-11, 3.88836e-11, 
    3.891827e-11, 3.898097e-11, 3.912475e-11, 3.904715e-11, 3.91379e-11, 
    3.893741e-11, 3.883333e-11, 3.880642e-11, 3.875616e-11, 3.880756e-11, 
    3.880338e-11, 3.885256e-11, 3.883676e-11, 3.895481e-11, 3.88914e-11, 
    3.90715e-11, 3.913719e-11, 3.932268e-11, 3.943634e-11, 3.955202e-11, 
    3.960308e-11, 3.961862e-11, 3.962512e-11 ;

 SOILC =
  17.34412, 17.34411, 17.34411, 17.3441, 17.34411, 17.3441, 17.34412, 
    17.34411, 17.34411, 17.34412, 17.34409, 17.3441, 17.34407, 17.34408, 
    17.34406, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34404, 
    17.34405, 17.34403, 17.34404, 17.34404, 17.34405, 17.3441, 17.34409, 
    17.3441, 17.3441, 17.3441, 17.34411, 17.34411, 17.34412, 17.34412, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34409, 
    17.34406, 17.34407, 17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 
    17.34406, 17.34406, 17.34406, 17.34408, 17.34408, 17.3441, 17.34411, 
    17.34412, 17.34412, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 
    17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34406, 17.34409, 17.3441, 17.34411, 17.34411, 17.34412, 17.34411, 
    17.34412, 17.34411, 17.34411, 17.34411, 17.3441, 17.3441, 17.34407, 
    17.34409, 17.34406, 17.34406, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34404, 17.34405, 17.34404, 17.34406, 17.34405, 17.34411, 
    17.34411, 17.34411, 17.34411, 17.34411, 17.34412, 17.34411, 17.34411, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34406, 17.34406, 17.34406, 17.34406, 17.34404, 17.34406, 
    17.34404, 17.34404, 17.34405, 17.34404, 17.34411, 17.34411, 17.34412, 
    17.34411, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 17.3441, 
    17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34406, 17.34404, 17.34404, 
    17.34404, 17.34404, 17.34411, 17.34411, 17.34411, 17.3441, 17.34411, 
    17.3441, 17.34409, 17.34408, 17.34408, 17.34407, 17.34408, 17.34408, 
    17.34407, 17.34408, 17.34406, 17.34408, 17.34405, 17.34407, 17.34405, 
    17.34406, 17.34405, 17.34405, 17.34404, 17.34403, 17.34404, 17.34403, 
    17.3441, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34407, 
    17.34407, 17.34407, 17.34406, 17.34408, 17.34407, 17.34409, 17.34409, 
    17.34409, 17.3441, 17.34407, 17.34409, 17.34406, 17.34407, 17.34405, 
    17.34406, 17.34404, 17.34403, 17.34402, 17.34401, 17.3441, 17.3441, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34407, 17.34407, 17.34406, 
    17.34406, 17.34407, 17.34406, 17.34409, 17.34407, 17.3441, 17.34409, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.344, 17.34402, 17.3441, 17.3441, 17.34408, 17.34409, 
    17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34407, 17.34406, 17.34408, 17.34408, 17.34408, 17.34408, 
    17.34407, 17.34407, 17.34407, 17.34406, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.34409, 17.34408, 17.34408, 17.34408, 17.34406, 17.34407, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34406, 
    17.34407, 17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34405, 17.34407, 17.34406, 17.34406, 17.34406, 17.34408, 
    17.34406, 17.34408, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34406, 17.34407, 17.34407, 17.34407, 17.34408, 17.34408, 
    17.34408, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34403, 
    17.34404, 17.34403, 17.34404, 17.34402, 17.34406, 17.34404, 17.34407, 
    17.34407, 17.34406, 17.34405, 17.34406, 17.34405, 17.34407, 17.34408, 
    17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34408, 17.34406, 
    17.34407, 17.34405, 17.34405, 17.34403, 17.34402, 17.34401, 17.344, 
    17.344, 17.344 ;

 SOILC_HR =
  7.623549e-08, 7.644416e-08, 7.640361e-08, 7.657187e-08, 7.647855e-08, 
    7.658871e-08, 7.627782e-08, 7.645243e-08, 7.634097e-08, 7.62543e-08, 
    7.689825e-08, 7.657938e-08, 7.722948e-08, 7.702619e-08, 7.75368e-08, 
    7.719783e-08, 7.760514e-08, 7.752706e-08, 7.776212e-08, 7.769479e-08, 
    7.79953e-08, 7.77932e-08, 7.815109e-08, 7.794706e-08, 7.797897e-08, 
    7.778652e-08, 7.664359e-08, 7.685854e-08, 7.663084e-08, 7.66615e-08, 
    7.664775e-08, 7.648046e-08, 7.639613e-08, 7.621956e-08, 7.625163e-08, 
    7.638132e-08, 7.667528e-08, 7.657553e-08, 7.682698e-08, 7.682131e-08, 
    7.710113e-08, 7.697498e-08, 7.744517e-08, 7.731157e-08, 7.76976e-08, 
    7.760053e-08, 7.769304e-08, 7.766499e-08, 7.76934e-08, 7.755104e-08, 
    7.761204e-08, 7.748676e-08, 7.69986e-08, 7.714208e-08, 7.671404e-08, 
    7.64565e-08, 7.628547e-08, 7.616406e-08, 7.618123e-08, 7.621394e-08, 
    7.638208e-08, 7.654015e-08, 7.666058e-08, 7.674113e-08, 7.682049e-08, 
    7.706056e-08, 7.718769e-08, 7.747217e-08, 7.742086e-08, 7.750779e-08, 
    7.759088e-08, 7.773031e-08, 7.770736e-08, 7.776877e-08, 7.750553e-08, 
    7.768048e-08, 7.739163e-08, 7.747064e-08, 7.684195e-08, 7.660245e-08, 
    7.650053e-08, 7.64114e-08, 7.619442e-08, 7.634426e-08, 7.62852e-08, 
    7.642574e-08, 7.651501e-08, 7.647086e-08, 7.674333e-08, 7.663741e-08, 
    7.719521e-08, 7.6955e-08, 7.758118e-08, 7.743139e-08, 7.761709e-08, 
    7.752234e-08, 7.768467e-08, 7.753858e-08, 7.779164e-08, 7.784672e-08, 
    7.780908e-08, 7.79537e-08, 7.753048e-08, 7.769302e-08, 7.646963e-08, 
    7.647682e-08, 7.651037e-08, 7.636287e-08, 7.635385e-08, 7.621868e-08, 
    7.633896e-08, 7.639017e-08, 7.652019e-08, 7.659708e-08, 7.667015e-08, 
    7.683081e-08, 7.701018e-08, 7.726096e-08, 7.744111e-08, 7.756182e-08, 
    7.748781e-08, 7.755315e-08, 7.74801e-08, 7.744587e-08, 7.782607e-08, 
    7.76126e-08, 7.79329e-08, 7.791519e-08, 7.777024e-08, 7.791719e-08, 
    7.648188e-08, 7.644044e-08, 7.629653e-08, 7.640916e-08, 7.620396e-08, 
    7.631881e-08, 7.638484e-08, 7.66396e-08, 7.669559e-08, 7.674747e-08, 
    7.684995e-08, 7.698143e-08, 7.721203e-08, 7.741262e-08, 7.759571e-08, 
    7.75823e-08, 7.758702e-08, 7.762791e-08, 7.752661e-08, 7.764454e-08, 
    7.766432e-08, 7.761258e-08, 7.791282e-08, 7.782705e-08, 7.791481e-08, 
    7.785898e-08, 7.645392e-08, 7.652364e-08, 7.648596e-08, 7.65568e-08, 
    7.650689e-08, 7.672879e-08, 7.679531e-08, 7.710651e-08, 7.697884e-08, 
    7.718206e-08, 7.699949e-08, 7.703184e-08, 7.718864e-08, 7.700937e-08, 
    7.740154e-08, 7.713565e-08, 7.762949e-08, 7.7364e-08, 7.764613e-08, 
    7.759493e-08, 7.767972e-08, 7.775563e-08, 7.785115e-08, 7.802734e-08, 
    7.798656e-08, 7.813389e-08, 7.662758e-08, 7.671798e-08, 7.671004e-08, 
    7.680465e-08, 7.687462e-08, 7.702625e-08, 7.726938e-08, 7.717797e-08, 
    7.73458e-08, 7.737948e-08, 7.712452e-08, 7.728104e-08, 7.67785e-08, 
    7.685969e-08, 7.681136e-08, 7.663471e-08, 7.7199e-08, 7.690944e-08, 
    7.744408e-08, 7.728728e-08, 7.774481e-08, 7.751729e-08, 7.79641e-08, 
    7.815497e-08, 7.833466e-08, 7.85445e-08, 7.676734e-08, 7.670592e-08, 
    7.681592e-08, 7.696804e-08, 7.710922e-08, 7.729684e-08, 7.731605e-08, 
    7.735118e-08, 7.744221e-08, 7.751873e-08, 7.736227e-08, 7.753791e-08, 
    7.687849e-08, 7.722414e-08, 7.668267e-08, 7.684573e-08, 7.695908e-08, 
    7.690938e-08, 7.716753e-08, 7.722835e-08, 7.747545e-08, 7.734774e-08, 
    7.810785e-08, 7.777165e-08, 7.87043e-08, 7.844376e-08, 7.668445e-08, 
    7.676714e-08, 7.705483e-08, 7.691796e-08, 7.730937e-08, 7.740568e-08, 
    7.748397e-08, 7.758402e-08, 7.759483e-08, 7.765411e-08, 7.755698e-08, 
    7.765028e-08, 7.729724e-08, 7.745503e-08, 7.702198e-08, 7.712739e-08, 
    7.70789e-08, 7.70257e-08, 7.718989e-08, 7.736472e-08, 7.73685e-08, 
    7.742454e-08, 7.758241e-08, 7.731096e-08, 7.815116e-08, 7.763233e-08, 
    7.68573e-08, 7.701648e-08, 7.703925e-08, 7.697759e-08, 7.739602e-08, 
    7.724444e-08, 7.765266e-08, 7.754237e-08, 7.772309e-08, 7.763329e-08, 
    7.762007e-08, 7.750472e-08, 7.743289e-08, 7.725138e-08, 7.710367e-08, 
    7.698654e-08, 7.701378e-08, 7.714245e-08, 7.737543e-08, 7.75958e-08, 
    7.754753e-08, 7.770936e-08, 7.7281e-08, 7.746063e-08, 7.73912e-08, 
    7.757223e-08, 7.717554e-08, 7.751326e-08, 7.708917e-08, 7.712637e-08, 
    7.724142e-08, 7.747279e-08, 7.752402e-08, 7.757865e-08, 7.754495e-08, 
    7.738135e-08, 7.735456e-08, 7.723864e-08, 7.720661e-08, 7.711827e-08, 
    7.704512e-08, 7.711195e-08, 7.718212e-08, 7.738143e-08, 7.756099e-08, 
    7.77567e-08, 7.780461e-08, 7.803313e-08, 7.784707e-08, 7.815405e-08, 
    7.7893e-08, 7.834487e-08, 7.753288e-08, 7.788538e-08, 7.724667e-08, 
    7.731551e-08, 7.743999e-08, 7.772545e-08, 7.757139e-08, 7.775158e-08, 
    7.735351e-08, 7.714686e-08, 7.709342e-08, 7.699366e-08, 7.709571e-08, 
    7.708741e-08, 7.718505e-08, 7.715368e-08, 7.738805e-08, 7.726216e-08, 
    7.761973e-08, 7.775017e-08, 7.811844e-08, 7.834409e-08, 7.857378e-08, 
    7.867516e-08, 7.8706e-08, 7.871891e-08 ;

 SOILC_LOSS =
  7.623549e-08, 7.644416e-08, 7.640361e-08, 7.657187e-08, 7.647855e-08, 
    7.658871e-08, 7.627782e-08, 7.645243e-08, 7.634097e-08, 7.62543e-08, 
    7.689825e-08, 7.657938e-08, 7.722948e-08, 7.702619e-08, 7.75368e-08, 
    7.719783e-08, 7.760514e-08, 7.752706e-08, 7.776212e-08, 7.769479e-08, 
    7.79953e-08, 7.77932e-08, 7.815109e-08, 7.794706e-08, 7.797897e-08, 
    7.778652e-08, 7.664359e-08, 7.685854e-08, 7.663084e-08, 7.66615e-08, 
    7.664775e-08, 7.648046e-08, 7.639613e-08, 7.621956e-08, 7.625163e-08, 
    7.638132e-08, 7.667528e-08, 7.657553e-08, 7.682698e-08, 7.682131e-08, 
    7.710113e-08, 7.697498e-08, 7.744517e-08, 7.731157e-08, 7.76976e-08, 
    7.760053e-08, 7.769304e-08, 7.766499e-08, 7.76934e-08, 7.755104e-08, 
    7.761204e-08, 7.748676e-08, 7.69986e-08, 7.714208e-08, 7.671404e-08, 
    7.64565e-08, 7.628547e-08, 7.616406e-08, 7.618123e-08, 7.621394e-08, 
    7.638208e-08, 7.654015e-08, 7.666058e-08, 7.674113e-08, 7.682049e-08, 
    7.706056e-08, 7.718769e-08, 7.747217e-08, 7.742086e-08, 7.750779e-08, 
    7.759088e-08, 7.773031e-08, 7.770736e-08, 7.776877e-08, 7.750553e-08, 
    7.768048e-08, 7.739163e-08, 7.747064e-08, 7.684195e-08, 7.660245e-08, 
    7.650053e-08, 7.64114e-08, 7.619442e-08, 7.634426e-08, 7.62852e-08, 
    7.642574e-08, 7.651501e-08, 7.647086e-08, 7.674333e-08, 7.663741e-08, 
    7.719521e-08, 7.6955e-08, 7.758118e-08, 7.743139e-08, 7.761709e-08, 
    7.752234e-08, 7.768467e-08, 7.753858e-08, 7.779164e-08, 7.784672e-08, 
    7.780908e-08, 7.79537e-08, 7.753048e-08, 7.769302e-08, 7.646963e-08, 
    7.647682e-08, 7.651037e-08, 7.636287e-08, 7.635385e-08, 7.621868e-08, 
    7.633896e-08, 7.639017e-08, 7.652019e-08, 7.659708e-08, 7.667015e-08, 
    7.683081e-08, 7.701018e-08, 7.726096e-08, 7.744111e-08, 7.756182e-08, 
    7.748781e-08, 7.755315e-08, 7.74801e-08, 7.744587e-08, 7.782607e-08, 
    7.76126e-08, 7.79329e-08, 7.791519e-08, 7.777024e-08, 7.791719e-08, 
    7.648188e-08, 7.644044e-08, 7.629653e-08, 7.640916e-08, 7.620396e-08, 
    7.631881e-08, 7.638484e-08, 7.66396e-08, 7.669559e-08, 7.674747e-08, 
    7.684995e-08, 7.698143e-08, 7.721203e-08, 7.741262e-08, 7.759571e-08, 
    7.75823e-08, 7.758702e-08, 7.762791e-08, 7.752661e-08, 7.764454e-08, 
    7.766432e-08, 7.761258e-08, 7.791282e-08, 7.782705e-08, 7.791481e-08, 
    7.785898e-08, 7.645392e-08, 7.652364e-08, 7.648596e-08, 7.65568e-08, 
    7.650689e-08, 7.672879e-08, 7.679531e-08, 7.710651e-08, 7.697884e-08, 
    7.718206e-08, 7.699949e-08, 7.703184e-08, 7.718864e-08, 7.700937e-08, 
    7.740154e-08, 7.713565e-08, 7.762949e-08, 7.7364e-08, 7.764613e-08, 
    7.759493e-08, 7.767972e-08, 7.775563e-08, 7.785115e-08, 7.802734e-08, 
    7.798656e-08, 7.813389e-08, 7.662758e-08, 7.671798e-08, 7.671004e-08, 
    7.680465e-08, 7.687462e-08, 7.702625e-08, 7.726938e-08, 7.717797e-08, 
    7.73458e-08, 7.737948e-08, 7.712452e-08, 7.728104e-08, 7.67785e-08, 
    7.685969e-08, 7.681136e-08, 7.663471e-08, 7.7199e-08, 7.690944e-08, 
    7.744408e-08, 7.728728e-08, 7.774481e-08, 7.751729e-08, 7.79641e-08, 
    7.815497e-08, 7.833466e-08, 7.85445e-08, 7.676734e-08, 7.670592e-08, 
    7.681592e-08, 7.696804e-08, 7.710922e-08, 7.729684e-08, 7.731605e-08, 
    7.735118e-08, 7.744221e-08, 7.751873e-08, 7.736227e-08, 7.753791e-08, 
    7.687849e-08, 7.722414e-08, 7.668267e-08, 7.684573e-08, 7.695908e-08, 
    7.690938e-08, 7.716753e-08, 7.722835e-08, 7.747545e-08, 7.734774e-08, 
    7.810785e-08, 7.777165e-08, 7.87043e-08, 7.844376e-08, 7.668445e-08, 
    7.676714e-08, 7.705483e-08, 7.691796e-08, 7.730937e-08, 7.740568e-08, 
    7.748397e-08, 7.758402e-08, 7.759483e-08, 7.765411e-08, 7.755698e-08, 
    7.765028e-08, 7.729724e-08, 7.745503e-08, 7.702198e-08, 7.712739e-08, 
    7.70789e-08, 7.70257e-08, 7.718989e-08, 7.736472e-08, 7.73685e-08, 
    7.742454e-08, 7.758241e-08, 7.731096e-08, 7.815116e-08, 7.763233e-08, 
    7.68573e-08, 7.701648e-08, 7.703925e-08, 7.697759e-08, 7.739602e-08, 
    7.724444e-08, 7.765266e-08, 7.754237e-08, 7.772309e-08, 7.763329e-08, 
    7.762007e-08, 7.750472e-08, 7.743289e-08, 7.725138e-08, 7.710367e-08, 
    7.698654e-08, 7.701378e-08, 7.714245e-08, 7.737543e-08, 7.75958e-08, 
    7.754753e-08, 7.770936e-08, 7.7281e-08, 7.746063e-08, 7.73912e-08, 
    7.757223e-08, 7.717554e-08, 7.751326e-08, 7.708917e-08, 7.712637e-08, 
    7.724142e-08, 7.747279e-08, 7.752402e-08, 7.757865e-08, 7.754495e-08, 
    7.738135e-08, 7.735456e-08, 7.723864e-08, 7.720661e-08, 7.711827e-08, 
    7.704512e-08, 7.711195e-08, 7.718212e-08, 7.738143e-08, 7.756099e-08, 
    7.77567e-08, 7.780461e-08, 7.803313e-08, 7.784707e-08, 7.815405e-08, 
    7.7893e-08, 7.834487e-08, 7.753288e-08, 7.788538e-08, 7.724667e-08, 
    7.731551e-08, 7.743999e-08, 7.772545e-08, 7.757139e-08, 7.775158e-08, 
    7.735351e-08, 7.714686e-08, 7.709342e-08, 7.699366e-08, 7.709571e-08, 
    7.708741e-08, 7.718505e-08, 7.715368e-08, 7.738805e-08, 7.726216e-08, 
    7.761973e-08, 7.775017e-08, 7.811844e-08, 7.834409e-08, 7.857378e-08, 
    7.867516e-08, 7.8706e-08, 7.871891e-08 ;

 SOILICE =
  98.96838, 99.4036, 99.31889, 99.67061, 99.47539, 99.70584, 99.0565, 
    99.42092, 99.18818, 99.00748, 100.3553, 99.68631, 101.0529, 100.6242, 
    101.703, 100.9861, 101.8479, 101.6823, 102.1812, 102.0381, 102.678, 
    102.2473, 103.0105, 102.575, 102.6431, 102.2331, 99.82069, 100.2719, 
    99.794, 99.85826, 99.82941, 99.47944, 99.30339, 98.93512, 99.00191, 
    99.2724, 99.88716, 99.67819, 100.2052, 100.1933, 100.782, 100.5163, 
    101.5088, 101.2261, 102.0441, 101.8381, 102.0344, 101.9749, 102.0352, 
    101.7331, 101.8625, 101.5968, 100.5661, 100.8684, 99.96835, 99.42953, 
    99.07247, 98.81961, 98.85533, 98.92347, 99.27399, 99.60417, 99.85625, 
    100.0251, 100.1916, 100.6968, 100.9647, 101.566, 101.4573, 101.6415, 
    101.8176, 102.1136, 102.0649, 102.1954, 101.6366, 102.0078, 101.3954, 
    101.5627, 100.2371, 99.73454, 99.52153, 99.33517, 98.88281, 99.19508, 
    99.07191, 99.36505, 99.55161, 99.4593, 100.0297, 99.80773, 100.9805, 
    100.4744, 101.797, 101.4796, 101.8732, 101.6722, 102.0167, 101.7066, 
    102.244, 102.3613, 102.2812, 102.5891, 101.6895, 102.0345, 99.45673, 
    99.47178, 99.54189, 99.2339, 99.21507, 98.9333, 99.18398, 99.29086, 
    99.56241, 99.72327, 99.87633, 100.2133, 100.5905, 101.1193, 101.5002, 
    101.7559, 101.599, 101.7375, 101.5827, 101.5102, 102.3174, 101.8637, 
    102.5448, 102.507, 102.1986, 102.5113, 99.48235, 99.39575, 99.09551, 
    99.33043, 98.90264, 99.14198, 99.27977, 99.81241, 99.92961, 100.0384, 
    100.2535, 100.5299, 101.0159, 101.4399, 101.8278, 101.7993, 101.8094, 
    101.8961, 101.6813, 101.9314, 101.9735, 101.8636, 102.502, 102.3194, 
    102.5062, 102.3873, 99.42389, 99.56964, 99.49087, 99.63903, 99.53465, 
    99.99934, 100.1389, 100.7935, 100.5245, 100.9527, 100.5679, 100.6361, 
    100.9668, 100.5887, 101.4165, 100.8549, 101.8995, 101.3372, 101.9348, 
    101.8261, 102.0061, 102.1675, 102.3707, 102.7463, 102.6592, 102.9737, 
    99.78714, 99.97663, 99.95991, 100.1584, 100.3054, 100.6243, 101.137, 
    100.944, 101.2985, 101.3697, 100.8313, 101.1617, 100.1035, 100.2741, 
    100.1725, 99.80209, 100.9885, 100.3786, 101.5065, 101.1748, 102.1445, 
    101.6616, 102.6113, 103.0189, 103.4032, 103.8535, 100.0801, 99.95125, 
    100.182, 100.5019, 100.7991, 101.195, 101.2356, 101.3099, 101.5025, 
    101.6646, 101.3334, 101.7052, 100.3137, 101.0415, 99.90259, 100.2448, 
    100.483, 100.3784, 100.922, 101.0503, 101.5729, 101.3026, 102.9183, 
    102.2016, 104.197, 103.6372, 99.90626, 100.0796, 100.6845, 100.3964, 
    101.2215, 101.4252, 101.5909, 101.8031, 101.826, 101.9518, 101.7456, 
    101.9436, 101.1959, 101.5296, 100.6152, 100.8374, 100.7351, 100.6231, 
    100.9691, 101.3386, 101.3465, 101.4651, 101.8001, 101.2248, 103.0111, 
    101.9059, 100.2689, 100.6038, 100.6517, 100.5218, 101.4047, 101.0843, 
    101.9487, 101.7147, 102.0983, 101.9076, 101.8795, 101.6349, 101.4828, 
    101.099, 100.7874, 100.5406, 100.598, 100.8691, 101.3613, 101.828, 
    101.7257, 102.0691, 101.1615, 101.5415, 101.3946, 101.778, 100.9389, 
    101.6534, 100.7568, 100.8352, 101.078, 101.5674, 101.6758, 101.7917, 
    101.7201, 101.3737, 101.317, 101.072, 101.0045, 100.8181, 100.6639, 
    100.8048, 100.9528, 101.3739, 101.7542, 102.1698, 102.2716, 102.7588, 
    102.3622, 103.0173, 102.4603, 103.4255, 101.6948, 102.4438, 101.089, 
    101.2344, 101.4979, 102.1035, 101.7762, 102.159, 101.3148, 100.8785, 
    100.7657, 100.5556, 100.7705, 100.7531, 100.9589, 100.8927, 101.3879, 
    101.1217, 101.8788, 102.1559, 102.9407, 103.4236, 103.9163, 104.1342, 
    104.2006, 104.2284,
  115.4026, 115.8126, 115.7328, 116.064, 115.8802, 116.0972, 115.4856, 
    115.829, 115.6097, 115.4395, 116.7084, 116.0788, 117.3639, 116.961, 
    117.9743, 117.3012, 118.1103, 117.9547, 118.4228, 118.2886, 118.8887, 
    118.4848, 119.2001, 118.7921, 118.8559, 118.4715, 116.2053, 116.63, 
    116.1801, 116.2406, 116.2135, 115.884, 115.7183, 115.3713, 115.4342, 
    115.6891, 116.2679, 116.0711, 116.567, 116.5558, 117.1093, 116.8596, 
    117.7919, 117.5265, 118.2942, 118.1009, 118.2852, 118.2293, 118.2859, 
    118.0024, 118.1238, 117.8746, 116.9064, 117.1905, 116.3442, 115.8372, 
    115.5007, 115.2624, 115.2961, 115.3603, 115.6906, 116.0014, 116.2387, 
    116.3976, 116.5542, 117.0294, 117.281, 117.8457, 117.7436, 117.9165, 
    118.0817, 118.3595, 118.3137, 118.4362, 117.9119, 118.2602, 117.6854, 
    117.8425, 116.5972, 116.1242, 115.9238, 115.7482, 115.322, 115.6162, 
    115.5002, 115.7763, 115.952, 115.865, 116.4019, 116.1931, 117.2959, 
    116.8202, 118.0624, 117.7645, 118.1339, 117.9453, 118.2685, 117.9776, 
    118.4817, 118.5917, 118.5166, 118.8052, 117.9615, 118.2852, 115.8626, 
    115.8768, 115.9428, 115.6528, 115.6351, 115.3696, 115.6058, 115.7064, 
    115.9621, 116.1136, 116.2576, 116.5747, 116.9294, 117.4262, 117.7838, 
    118.0238, 117.8766, 118.0066, 117.8613, 117.7932, 118.5505, 118.125, 
    118.7637, 118.7283, 118.4391, 118.7323, 115.8867, 115.8052, 115.5224, 
    115.7437, 115.3407, 115.5662, 115.696, 116.1975, 116.3077, 116.4101, 
    116.6124, 116.8724, 117.3291, 117.7273, 118.0913, 118.0646, 118.074, 
    118.1554, 117.9538, 118.1885, 118.228, 118.1249, 118.7235, 118.5524, 
    118.7275, 118.616, 115.8317, 115.9689, 115.8948, 116.0343, 115.936, 
    116.3734, 116.5047, 117.1202, 116.8673, 117.2698, 116.9081, 116.9722, 
    117.2831, 116.9276, 117.7054, 117.1779, 118.1586, 117.631, 118.1917, 
    118.0897, 118.2586, 118.41, 118.6005, 118.9525, 118.8709, 119.1656, 
    116.1737, 116.352, 116.3362, 116.523, 116.6612, 116.961, 117.4428, 
    117.2615, 117.5944, 117.6614, 117.1556, 117.466, 116.4714, 116.6319, 
    116.5363, 116.1878, 117.3034, 116.7302, 117.7897, 117.4783, 118.3884, 
    117.9354, 118.826, 119.2081, 119.5678, 119.9893, 116.4493, 116.3281, 
    116.5452, 116.846, 117.1253, 117.4973, 117.5354, 117.6052, 117.786, 
    117.9381, 117.6273, 117.9763, 116.6693, 117.3532, 116.2823, 116.6043, 
    116.8283, 116.7299, 117.2408, 117.3614, 117.8522, 117.5983, 119.1138, 
    118.4421, 120.3105, 119.7869, 116.2858, 116.4489, 117.0177, 116.7469, 
    117.5221, 117.7134, 117.869, 118.0681, 118.0896, 118.2076, 118.0142, 
    118.2, 117.4981, 117.8115, 116.9525, 117.1613, 117.0652, 116.9599, 
    117.2851, 117.6322, 117.6395, 117.751, 118.0656, 117.5253, 119.2009, 
    118.1648, 116.6269, 116.9419, 116.9868, 116.8647, 117.6942, 117.3933, 
    118.2047, 117.9851, 118.345, 118.1661, 118.1398, 117.9102, 117.7675, 
    117.4071, 117.1144, 116.8824, 116.9363, 117.1912, 117.6535, 118.0916, 
    117.9955, 118.3176, 117.4658, 117.8227, 117.6847, 118.0446, 117.2567, 
    117.9279, 117.0855, 117.1592, 117.3874, 117.847, 117.9486, 118.0574, 
    117.9903, 117.6652, 117.6119, 117.3818, 117.3184, 117.1432, 116.9983, 
    117.1307, 117.2698, 117.6653, 118.0223, 118.4121, 118.5076, 118.9644, 
    118.5927, 119.2067, 118.6848, 119.5888, 117.9666, 118.6692, 117.3977, 
    117.5343, 117.7817, 118.35, 118.0429, 118.402, 117.6098, 117.2, 117.094, 
    116.8965, 117.0985, 117.0821, 117.2755, 117.2133, 117.6784, 117.4285, 
    118.1392, 118.3992, 119.1348, 119.5869, 120.0479, 120.2518, 120.3138, 
    120.3398,
  168.5735, 169.1529, 169.0401, 169.5082, 169.2484, 169.5551, 168.6908, 
    169.176, 168.8661, 168.6255, 170.419, 169.5291, 171.3455, 170.776, 
    172.2084, 171.2569, 172.4006, 172.1807, 172.8425, 172.6527, 173.501, 
    172.9301, 173.9414, 173.3645, 173.4547, 172.9113, 169.7078, 170.3081, 
    169.6723, 169.7578, 169.7194, 169.2538, 169.0196, 168.5291, 168.6181, 
    168.9783, 169.7963, 169.5182, 170.2192, 170.2033, 170.9857, 170.6327, 
    171.9505, 171.5753, 172.6606, 172.3874, 172.6478, 172.5688, 172.6488, 
    172.2482, 172.4198, 172.0674, 170.6988, 171.1004, 169.9042, 169.1875, 
    168.7121, 168.3753, 168.4229, 168.5136, 168.9804, 169.4198, 169.7551, 
    169.9796, 170.201, 170.8726, 171.2283, 172.0265, 171.8822, 172.1266, 
    172.3602, 172.7529, 172.6882, 172.8613, 172.1201, 172.6126, 171.8, 
    172.0221, 170.2618, 169.5932, 169.31, 169.0618, 168.4595, 168.8753, 
    168.7113, 169.1015, 169.3498, 169.227, 169.9858, 169.6906, 171.2494, 
    170.577, 172.3329, 171.9118, 172.4339, 172.1674, 172.6243, 172.213, 
    172.9257, 173.0812, 172.975, 173.3831, 172.1903, 172.6479, 169.2236, 
    169.2436, 169.3369, 168.927, 168.9019, 168.5267, 168.8605, 169.0028, 
    169.3642, 169.5782, 169.7818, 170.2299, 170.7313, 171.4336, 171.9391, 
    172.2784, 172.0703, 172.254, 172.0486, 171.9524, 173.023, 172.4214, 
    173.3244, 173.2743, 172.8654, 173.2799, 169.2577, 169.1424, 168.7427, 
    169.0555, 168.4859, 168.8046, 168.9881, 169.6969, 169.8527, 169.9974, 
    170.2833, 170.6507, 171.2964, 171.8592, 172.3737, 172.336, 172.3493, 
    172.4644, 172.1794, 172.5112, 172.567, 172.4213, 173.2676, 173.0256, 
    173.2732, 173.1156, 169.1798, 169.3738, 169.269, 169.4662, 169.3273, 
    169.9455, 170.1311, 171.001, 170.6435, 171.2124, 170.7012, 170.7918, 
    171.2312, 170.7288, 171.8282, 171.0826, 172.4689, 171.723, 172.5157, 
    172.3715, 172.6102, 172.8242, 173.0936, 173.5913, 173.476, 173.8926, 
    169.6632, 169.9153, 169.893, 170.1569, 170.3523, 170.776, 171.4571, 
    171.2008, 171.6714, 171.766, 171.051, 171.4899, 170.084, 170.3108, 
    170.1757, 169.6831, 171.26, 170.4497, 171.9475, 171.5072, 172.7937, 
    172.1534, 173.4125, 173.9526, 174.4613, 175.0573, 170.0528, 169.8814, 
    170.1883, 170.6135, 171.0083, 171.5341, 171.5879, 171.6866, 171.9421, 
    172.1572, 171.7179, 172.2112, 170.3636, 171.3303, 169.8168, 170.2719, 
    170.5884, 170.4494, 171.1715, 171.3419, 172.0357, 171.6768, 173.8193, 
    172.8696, 175.5115, 174.7711, 169.8216, 170.0522, 170.8562, 170.4733, 
    171.5692, 171.8396, 172.0595, 172.341, 172.3713, 172.5382, 172.2648, 
    172.5274, 171.5352, 171.9782, 170.764, 171.0592, 170.9233, 170.7745, 
    171.2341, 171.7248, 171.7351, 171.8927, 172.3373, 171.5736, 173.9424, 
    172.4777, 170.3038, 170.749, 170.8125, 170.6399, 171.8125, 171.3871, 
    172.5341, 172.2237, 172.7325, 172.4795, 172.4424, 172.1178, 171.916, 
    171.4066, 170.9928, 170.6649, 170.7411, 171.1013, 171.7548, 172.3741, 
    172.2384, 172.6938, 171.4896, 171.994, 171.799, 172.3077, 171.194, 
    172.1427, 170.9521, 171.0562, 171.3787, 172.0284, 172.1721, 172.3259, 
    172.2309, 171.7714, 171.6961, 171.3708, 171.2811, 171.0335, 170.8288, 
    171.0159, 171.2125, 171.7715, 172.2762, 172.8273, 172.9623, 173.6082, 
    173.0825, 173.9506, 173.2128, 174.491, 172.1975, 173.1908, 171.3933, 
    171.5864, 171.9361, 172.7395, 172.3053, 172.813, 171.6931, 171.1139, 
    170.964, 170.6849, 170.9704, 170.9471, 171.2206, 171.1327, 171.7901, 
    171.4368, 172.4415, 172.809, 173.849, 174.4883, 175.1402, 175.4285, 
    175.5162, 175.5529,
  257.5481, 258.4214, 258.2544, 258.9476, 258.5629, 259.0171, 257.7278, 
    258.4556, 257.9964, 257.6278, 260.2971, 258.9786, 261.6711, 260.8264, 
    262.9517, 261.5396, 263.2371, 262.9107, 263.8934, 263.6116, 264.872, 
    264.0236, 265.5267, 264.6691, 264.8032, 263.9957, 259.2433, 260.1327, 
    259.1907, 259.3174, 259.2605, 258.5709, 258.224, 257.4802, 257.6165, 
    258.1628, 259.3744, 258.9625, 260.001, 259.9775, 261.1374, 260.614, 
    262.569, 262.0122, 263.6234, 263.2175, 263.6043, 263.487, 263.6059, 
    263.0108, 263.2657, 262.7424, 260.712, 261.3076, 259.5343, 258.4726, 
    257.7604, 257.2446, 257.3175, 257.4565, 258.166, 258.8167, 259.3134, 
    259.6461, 259.9742, 260.9697, 261.4973, 262.6818, 262.4676, 262.8304, 
    263.1772, 263.7603, 263.6642, 263.9214, 262.8207, 263.5519, 262.3456, 
    262.6752, 260.0641, 259.0735, 258.6539, 258.2865, 257.3735, 258.0104, 
    257.7593, 258.3454, 258.713, 258.5311, 259.6552, 259.2178, 261.5286, 
    260.5314, 263.1367, 262.5115, 263.2867, 262.8909, 263.5694, 262.9587, 
    264.0172, 264.2481, 264.0903, 264.6967, 262.9249, 263.6044, 258.5261, 
    258.5557, 258.6939, 258.0869, 258.0498, 257.4765, 257.9878, 258.1992, 
    258.7343, 259.0514, 259.353, 260.017, 260.7602, 261.8019, 262.552, 
    263.0558, 262.7467, 263.0196, 262.7146, 262.5717, 264.1616, 263.2681, 
    264.6095, 264.5351, 263.9276, 264.5435, 258.5766, 258.4059, 257.8074, 
    258.2771, 257.414, 257.9022, 258.1774, 259.2271, 259.4579, 259.6724, 
    260.0961, 260.6408, 261.5983, 262.4334, 263.1973, 263.1413, 263.161, 
    263.332, 262.9088, 263.4015, 263.4843, 263.2679, 264.5251, 264.1655, 
    264.5335, 264.2993, 258.4613, 258.7486, 258.5934, 258.8853, 258.6797, 
    259.5954, 259.8705, 261.1601, 260.6301, 261.4738, 260.7156, 260.8499, 
    261.5016, 260.7565, 262.3874, 261.2811, 263.3386, 262.2312, 263.4081, 
    263.194, 263.5485, 263.8664, 264.2665, 265.0062, 264.8348, 265.4542, 
    259.1772, 259.5507, 259.5176, 259.9088, 260.1983, 260.8266, 261.8367, 
    261.4565, 262.1547, 262.2951, 261.2344, 261.8854, 259.8007, 260.1368, 
    259.9366, 259.2067, 261.5443, 260.3428, 262.5645, 261.9112, 263.821, 
    262.8701, 264.7405, 265.5433, 266.3, 267.1869, 259.7545, 259.5006, 
    259.9553, 260.5855, 261.171, 261.951, 262.0308, 262.1772, 262.5565, 
    262.8758, 262.2237, 262.9559, 260.2151, 261.6487, 259.4047, 260.0791, 
    260.5483, 260.3423, 261.413, 261.6659, 262.6954, 262.1628, 265.3451, 
    263.9337, 267.8632, 266.7609, 259.4119, 259.7536, 260.9454, 260.3778, 
    262.0031, 262.4043, 262.7307, 263.1487, 263.1937, 263.4416, 263.0355, 
    263.4254, 261.9527, 262.61, 260.8088, 261.2464, 261.045, 260.8242, 
    261.506, 262.2339, 262.2493, 262.4831, 263.1431, 262.0096, 265.5281, 
    263.3515, 260.1265, 260.7865, 260.8806, 260.6248, 262.3641, 261.7329, 
    263.4355, 262.9745, 263.7301, 263.3544, 263.2992, 262.8174, 262.5177, 
    261.7619, 261.148, 260.6618, 260.7748, 261.309, 262.2785, 263.1979, 
    262.9963, 263.6726, 261.885, 262.6336, 262.3441, 263.0993, 261.4464, 
    262.8541, 261.0876, 261.2421, 261.7204, 262.6845, 262.8979, 263.1262, 
    262.9853, 262.3031, 262.1913, 261.7087, 261.5757, 261.2084, 260.9048, 
    261.1823, 261.4739, 262.3033, 263.0524, 263.8709, 264.0714, 265.0312, 
    264.25, 265.5403, 264.4434, 266.344, 262.9355, 264.4108, 261.7421, 
    262.0286, 262.5476, 263.7404, 263.0958, 263.8497, 262.187, 261.3275, 
    261.1053, 260.6914, 261.1148, 261.0803, 261.4859, 261.3555, 262.3308, 
    261.8066, 263.2979, 263.8437, 265.3893, 266.3401, 267.3103, 267.7395, 
    267.8702, 267.9249,
  404.2867, 405.7206, 405.4413, 406.6009, 405.9572, 406.7171, 404.5769, 
    405.7776, 405.0107, 404.4155, 408.8613, 406.6527, 411.1056, 409.7352, 
    413.1868, 410.8921, 413.6511, 413.1202, 414.7199, 414.2609, 416.3148, 
    414.9319, 417.3835, 415.9839, 416.2026, 414.8864, 407.096, 408.5857, 
    407.0079, 407.22, 407.1248, 405.9706, 405.3903, 404.1772, 404.3972, 
    405.2882, 407.3153, 406.6259, 408.3654, 408.326, 410.2396, 409.3907, 
    412.5645, 411.6598, 414.2801, 413.6194, 414.249, 414.058, 414.2515, 
    413.2831, 413.6977, 412.8466, 409.5496, 410.5157, 407.5833, 405.806, 
    404.6295, 403.797, 403.9146, 404.1389, 405.2934, 406.3818, 407.2133, 
    407.7706, 408.3203, 409.9673, 410.8235, 412.7479, 412.3997, 412.9896, 
    413.5537, 414.503, 414.3466, 414.7654, 412.9739, 414.1637, 412.2015, 
    412.7372, 408.4706, 406.8117, 406.1093, 405.495, 404.005, 405.0334, 
    404.6277, 405.5935, 406.2085, 405.9041, 407.7858, 407.0532, 410.8743, 
    409.2545, 413.4879, 412.4711, 413.732, 413.088, 414.1921, 413.1983, 
    414.9214, 415.2977, 415.0405, 416.0291, 413.1433, 414.2491, 405.8957, 
    405.9453, 406.1765, 405.1613, 405.0993, 404.1713, 404.9968, 405.349, 
    406.2441, 406.7746, 407.2796, 408.3921, 409.6277, 411.3181, 412.537, 
    413.3562, 412.8536, 413.2973, 412.8014, 412.5691, 415.1567, 413.7016, 
    415.8868, 415.7655, 414.7755, 415.7792, 405.9801, 405.6947, 404.7054, 
    405.4794, 404.0703, 404.8585, 405.3125, 407.0687, 407.4554, 407.8146, 
    408.5247, 409.4341, 410.9875, 412.3441, 413.5865, 413.4954, 413.5275, 
    413.8056, 413.1171, 413.9188, 414.0536, 413.7014, 415.7493, 415.1631, 
    415.763, 415.3811, 405.7874, 406.2679, 406.0082, 406.4968, 406.1526, 
    407.6856, 408.1464, 410.2762, 409.4168, 410.7853, 409.5555, 409.7732, 
    410.8304, 409.6219, 412.2693, 410.4727, 413.8165, 412.0154, 413.9296, 
    413.5812, 414.1582, 414.6758, 415.3278, 416.5339, 416.2543, 417.265, 
    406.9853, 407.6106, 407.5554, 408.2107, 408.696, 409.7355, 411.3747, 
    410.7574, 411.8913, 412.1194, 410.3969, 411.4537, 408.0296, 408.5928, 
    408.2573, 407.0346, 410.8997, 408.9381, 412.5572, 411.4956, 414.6019, 
    413.0541, 416.1004, 417.4105, 418.6469, 420.0977, 407.9522, 407.5268, 
    408.2886, 409.3445, 410.294, 411.5603, 411.69, 411.9278, 412.5443, 
    413.0635, 412.0032, 413.1938, 408.7238, 411.0693, 407.3662, 408.4961, 
    409.2829, 408.9374, 410.6869, 411.0974, 412.7701, 411.9044, 417.0869, 
    414.7854, 421.2055, 419.4006, 407.3783, 407.9507, 409.928, 408.997, 
    411.6449, 412.2969, 412.8276, 413.5073, 413.5806, 413.984, 413.3233, 
    413.9578, 411.563, 412.6313, 409.7066, 410.4165, 410.0897, 409.7317, 
    410.8377, 412.0199, 412.045, 412.4249, 413.4978, 411.6556, 417.3853, 
    413.8371, 408.5757, 409.6703, 409.823, 409.4082, 412.2315, 411.2061, 
    413.9741, 413.224, 414.4538, 413.8422, 413.7523, 412.9684, 412.4812, 
    411.2531, 410.2567, 409.4683, 409.6515, 410.518, 412.0923, 413.5874, 
    413.2594, 414.3602, 411.4531, 412.6695, 412.199, 413.427, 410.7411, 
    413.0278, 410.1588, 410.4095, 411.1858, 412.7523, 413.0994, 413.4708, 
    413.2415, 412.1323, 411.9507, 411.1668, 410.9508, 410.3549, 409.8623, 
    410.3123, 410.7856, 412.1327, 413.3507, 414.6832, 415.0099, 416.5744, 
    415.3006, 417.4052, 415.6156, 418.7186, 413.1604, 415.5627, 411.2211, 
    411.6864, 412.5297, 414.4705, 413.4213, 414.6485, 411.9436, 410.548, 
    410.1875, 409.5163, 410.2029, 410.147, 410.8051, 410.5935, 412.1775, 
    411.3258, 413.7501, 414.6387, 417.1591, 418.7125, 420.2999, 421.0029, 
    421.2171, 421.3067,
  676.3514, 678.8893, 678.3947, 680.4435, 679.3086, 680.6429, 676.8647, 
    678.9904, 677.6322, 676.5792, 684.3256, 680.5323, 688.2996, 685.8549, 
    692.0219, 687.9184, 692.8539, 691.9026, 694.7712, 693.9474, 697.6378, 
    695.1519, 699.5627, 697.0427, 697.4361, 695.0702, 681.2928, 683.8516, 
    681.1418, 681.5056, 681.3423, 679.3322, 678.3042, 676.1578, 676.5467, 
    678.1234, 681.6693, 680.4865, 683.4731, 683.4055, 686.7542, 685.2411, 
    690.9078, 689.2897, 693.9818, 692.7971, 693.9261, 693.5834, 693.9306, 
    692.1944, 692.9374, 691.4127, 685.5242, 687.2466, 682.1293, 679.0406, 
    676.9578, 675.4857, 675.6935, 676.09, 678.1327, 680.0613, 681.4943, 
    682.451, 683.3957, 686.2684, 687.7959, 691.2359, 690.6129, 691.6687, 
    692.6794, 694.3819, 694.1012, 694.853, 691.6406, 693.773, 690.2584, 
    691.2169, 683.6538, 680.8052, 679.5782, 678.4897, 675.8533, 677.6724, 
    676.9545, 678.6642, 679.754, 679.2146, 682.4772, 681.2195, 687.8866, 
    685.0024, 692.5614, 690.7407, 692.9989, 691.8451, 693.824, 692.0426, 
    695.133, 695.809, 695.3469, 697.1241, 691.9441, 693.9262, 679.1996, 
    679.2875, 679.6973, 677.8989, 677.789, 676.1472, 677.6077, 678.2311, 
    679.8172, 680.7415, 681.608, 683.519, 685.6633, 688.6791, 690.8585, 
    692.3255, 691.4253, 692.2199, 691.3317, 690.916, 695.5556, 692.9445, 
    696.868, 696.65, 694.8709, 696.6745, 679.3492, 678.8434, 677.092, 
    678.4621, 675.9688, 677.3629, 678.1664, 681.246, 681.9099, 682.5266, 
    683.7471, 685.3185, 688.0887, 690.5133, 692.7382, 692.5748, 692.6324, 
    693.1309, 691.8971, 693.3338, 693.5755, 692.944, 696.6207, 695.5671, 
    696.6453, 695.959, 679.0078, 679.8594, 679.399, 680.265, 679.6549, 
    682.305, 683.0966, 686.8195, 685.2875, 687.7278, 685.5347, 685.9226, 
    687.8081, 685.6529, 690.3795, 687.1698, 693.1503, 689.9252, 693.3532, 
    692.7286, 693.7632, 694.692, 695.863, 698.0324, 697.5291, 699.3493, 
    681.103, 682.1763, 682.0815, 683.2072, 684.0416, 685.8553, 688.7803, 
    687.6781, 689.7036, 690.1114, 687.0349, 688.9214, 682.8959, 683.8641, 
    683.2872, 681.1876, 687.9321, 684.458, 690.8946, 688.9964, 694.5594, 
    691.7842, 697.2523, 699.6114, 701.8425, 704.4656, 682.763, 682.0324, 
    683.3412, 685.1587, 686.8513, 689.112, 689.3438, 689.7689, 690.8717, 
    691.8012, 689.9036, 692.0345, 684.0892, 688.2349, 681.7567, 683.6976, 
    685.0513, 684.4568, 687.5522, 688.285, 691.2756, 689.7271, 699.0281, 
    694.8886, 706.4728, 703.2045, 681.7775, 682.7604, 686.1985, 684.5593, 
    689.2632, 690.429, 691.3787, 692.5961, 692.7276, 693.4507, 692.2664, 
    693.4038, 689.1168, 691.0273, 685.804, 687.0697, 686.4869, 685.8487, 
    687.8215, 689.9335, 689.9784, 690.6579, 692.5788, 689.2823, 699.5658, 
    693.187, 683.8347, 685.7391, 686.0114, 685.2723, 690.312, 688.4792, 
    693.433, 692.0886, 694.2935, 693.1965, 693.0353, 691.6309, 690.7588, 
    688.5632, 686.7847, 685.3794, 685.7057, 687.2509, 690.0629, 692.7397, 
    692.1519, 694.1255, 688.9205, 691.0957, 690.2538, 692.4524, 687.6489, 
    691.7369, 686.6102, 687.0572, 688.4429, 691.2438, 691.8655, 692.5307, 
    692.1201, 690.1345, 689.8099, 688.4091, 688.0233, 686.9598, 686.0814, 
    686.884, 687.7285, 690.1352, 692.3156, 694.7052, 695.2919, 698.1051, 
    695.8141, 699.6016, 696.38, 701.9717, 691.9745, 696.285, 688.506, 
    689.3373, 690.8454, 694.3234, 692.442, 694.6429, 689.7972, 687.3044, 
    686.6614, 685.4648, 686.6888, 686.5891, 687.7632, 687.3856, 690.2153, 
    688.693, 693.0314, 694.6254, 699.1583, 701.9608, 704.8318, 706.1055, 
    706.4939, 706.6564,
  1152.656, 1157.944, 1156.912, 1161.209, 1158.821, 1161.641, 1153.723, 
    1158.156, 1155.322, 1153.129, 1169.655, 1161.402, 1178.195, 1172.999, 
    1186.158, 1177.383, 1187.946, 1185.902, 1192.08, 1190.302, 1198.293, 
    1192.903, 1202.487, 1197, 1197.854, 1192.726, 1163.052, 1168.62, 
    1162.724, 1163.513, 1163.159, 1158.87, 1156.723, 1152.254, 1153.062, 
    1156.346, 1163.869, 1161.302, 1167.795, 1167.647, 1174.907, 1171.657, 
    1183.768, 1180.307, 1190.376, 1187.824, 1190.256, 1189.517, 1190.266, 
    1186.529, 1188.126, 1184.85, 1172.276, 1175.954, 1164.869, 1158.261, 
    1153.917, 1150.858, 1151.289, 1152.113, 1156.365, 1160.396, 1163.489, 
    1165.569, 1167.626, 1173.876, 1177.122, 1184.471, 1183.136, 1185.4, 
    1187.571, 1191.24, 1190.634, 1192.257, 1185.339, 1189.926, 1182.378, 
    1184.431, 1168.189, 1161.993, 1159.384, 1157.11, 1151.621, 1155.406, 
    1153.91, 1157.474, 1159.752, 1158.624, 1165.626, 1162.892, 1177.316, 
    1171.135, 1187.317, 1183.41, 1188.259, 1185.778, 1190.036, 1186.203, 
    1192.862, 1194.325, 1193.325, 1197.177, 1185.991, 1190.256, 1158.593, 
    1158.777, 1159.634, 1155.877, 1155.648, 1152.231, 1155.271, 1156.571, 
    1159.885, 1161.855, 1163.736, 1167.895, 1172.581, 1179.004, 1183.662, 
    1186.81, 1184.877, 1186.583, 1184.677, 1183.786, 1193.776, 1188.141, 
    1196.621, 1196.147, 1192.296, 1196.201, 1158.906, 1157.849, 1154.197, 
    1157.052, 1151.861, 1154.76, 1156.436, 1162.95, 1164.392, 1165.733, 
    1168.392, 1171.826, 1177.746, 1182.923, 1187.698, 1187.346, 1187.47, 
    1188.543, 1185.89, 1188.98, 1189.5, 1188.14, 1196.084, 1193.801, 
    1196.137, 1194.65, 1158.192, 1159.973, 1159.01, 1160.823, 1159.545, 
    1165.251, 1166.974, 1175.046, 1171.758, 1176.978, 1172.299, 1173.143, 
    1177.148, 1172.558, 1182.637, 1175.791, 1188.584, 1181.665, 1189.021, 
    1187.677, 1189.905, 1191.909, 1194.442, 1199.151, 1198.056, 1202.021, 
    1162.639, 1164.971, 1164.765, 1167.215, 1169.035, 1173, 1179.22, 
    1176.872, 1181.191, 1182.063, 1175.504, 1179.521, 1166.537, 1168.648, 
    1167.39, 1162.823, 1177.412, 1169.944, 1183.74, 1179.681, 1191.623, 
    1185.648, 1197.455, 1202.593, 1207.477, 1213.251, 1166.248, 1164.658, 
    1167.507, 1171.476, 1175.114, 1179.928, 1180.423, 1181.331, 1183.691, 
    1185.684, 1181.619, 1186.185, 1169.139, 1178.057, 1164.059, 1168.285, 
    1171.241, 1169.942, 1176.604, 1178.164, 1184.557, 1181.241, 1201.32, 
    1192.334, 1217.694, 1210.471, 1164.104, 1166.242, 1173.728, 1170.166, 
    1180.251, 1182.743, 1184.778, 1187.392, 1187.675, 1189.231, 1186.683, 
    1189.13, 1179.938, 1184.024, 1172.889, 1175.578, 1174.34, 1172.986, 
    1177.177, 1181.683, 1181.779, 1183.233, 1187.355, 1180.292, 1202.493, 
    1188.663, 1168.583, 1172.747, 1173.331, 1171.725, 1182.492, 1178.578, 
    1189.193, 1186.301, 1191.049, 1188.684, 1188.337, 1185.318, 1183.449, 
    1178.757, 1174.972, 1171.959, 1172.674, 1175.963, 1181.959, 1187.701, 
    1186.437, 1190.686, 1179.519, 1184.171, 1182.368, 1187.083, 1176.81, 
    1185.546, 1174.602, 1175.551, 1178.501, 1184.488, 1185.822, 1187.251, 
    1186.369, 1182.113, 1181.418, 1178.429, 1177.607, 1175.344, 1173.48, 
    1175.183, 1176.979, 1182.114, 1186.789, 1191.938, 1193.206, 1199.309, 
    1194.336, 1202.572, 1195.562, 1207.761, 1186.056, 1195.356, 1178.635, 
    1180.409, 1183.635, 1191.113, 1187.061, 1191.803, 1181.391, 1176.077, 
    1174.71, 1172.146, 1174.769, 1174.557, 1177.053, 1176.25, 1182.286, 
    1179.034, 1188.328, 1191.765, 1201.604, 1207.737, 1214.061, 1216.879, 
    1217.741, 1218.101,
  2105.699, 2120.385, 2117.5, 2129.56, 2122.839, 2130.781, 2108.646, 
    2120.976, 2113.075, 2107.005, 2153.699, 2130.104, 2179.253, 2163.429, 
    2204.022, 2176.763, 2209.558, 2203.216, 2222.352, 2216.827, 2241.925, 
    2224.92, 2255.381, 2237.816, 2240.529, 2224.368, 2134.775, 2150.71, 
    2133.845, 2136.087, 2135.08, 2122.978, 2116.974, 2104.591, 2106.819, 
    2115.923, 2137.098, 2129.823, 2148.331, 2147.907, 2169.21, 2159.509, 
    2196.521, 2185.76, 2217.056, 2209.183, 2216.684, 2214.399, 2216.714, 
    2205.191, 2210.111, 2199.911, 2161.314, 2172.396, 2139.947, 2121.27, 
    2109.182, 2100.754, 2101.938, 2104.203, 2115.977, 2127.265, 2136.017, 
    2141.945, 2147.846, 2166.082, 2175.965, 2198.722, 2194.547, 2201.636, 
    2208.406, 2219.735, 2217.855, 2222.903, 2201.447, 2215.662, 2192.183, 
    2198.594, 2149.466, 2131.776, 2124.421, 2118.054, 2102.85, 2113.308, 
    2109.163, 2119.071, 2125.455, 2122.289, 2142.108, 2134.323, 2176.556, 
    2157.99, 2207.627, 2195.402, 2210.518, 2202.827, 2216.003, 2204.162, 
    2224.792, 2229.375, 2226.239, 2238.376, 2203.496, 2216.685, 2122.2, 
    2122.716, 2125.121, 2114.62, 2113.983, 2104.53, 2112.933, 2116.549, 
    2125.827, 2131.386, 2136.719, 2148.619, 2162.203, 2181.74, 2196.19, 
    2206.073, 2199.995, 2205.364, 2199.366, 2196.575, 2227.654, 2210.157, 
    2236.615, 2235.118, 2223.023, 2235.286, 2123.078, 2120.117, 2109.955, 
    2117.893, 2103.51, 2111.518, 2116.173, 2134.486, 2138.586, 2142.416, 
    2150.052, 2160.001, 2177.875, 2193.883, 2208.794, 2207.716, 2208.095, 
    2211.393, 2203.178, 2212.739, 2214.346, 2210.155, 2234.917, 2227.732, 
    2235.086, 2230.396, 2121.078, 2126.075, 2123.37, 2128.469, 2124.872, 
    2141.037, 2145.972, 2169.632, 2159.804, 2175.522, 2161.381, 2163.862, 
    2176.044, 2162.136, 2192.99, 2171.898, 2211.521, 2189.968, 2212.868, 
    2208.73, 2215.597, 2221.818, 2229.742, 2244.662, 2241.172, 2253.877, 
    2133.606, 2140.238, 2139.65, 2146.664, 2151.907, 2163.432, 2182.406, 
    2175.198, 2188.498, 2191.205, 2171.024, 2183.333, 2144.718, 2150.788, 
    2147.166, 2134.127, 2176.853, 2154.537, 2196.432, 2183.827, 2220.927, 
    2202.415, 2239.26, 2255.725, 2271.663, 2290.879, 2143.889, 2139.346, 
    2147.504, 2158.984, 2169.838, 2184.588, 2186.118, 2188.931, 2196.279, 
    2202.53, 2189.824, 2204.108, 2152.207, 2178.83, 2137.638, 2149.741, 
    2158.3, 2154.529, 2174.379, 2179.158, 2198.989, 2188.653, 2251.618, 
    2223.143, 2305.953, 2281.574, 2137.767, 2143.872, 2165.633, 2155.178, 
    2185.585, 2193.32, 2199.682, 2207.856, 2208.724, 2213.516, 2205.679, 
    2213.204, 2184.62, 2197.322, 2163.103, 2171.25, 2167.487, 2163.389, 
    2176.132, 2190.022, 2190.321, 2194.848, 2207.741, 2185.712, 2255.403, 
    2211.764, 2150.603, 2162.687, 2164.432, 2159.707, 2192.54, 2180.429, 
    2213.398, 2204.474, 2219.143, 2211.827, 2210.759, 2201.38, 2195.523, 
    2180.98, 2169.407, 2160.39, 2162.474, 2172.423, 2190.882, 2208.803, 
    2204.903, 2218.018, 2183.327, 2197.78, 2192.152, 2206.908, 2175.008, 
    2202.095, 2168.281, 2171.169, 2180.192, 2198.775, 2202.964, 2207.425, 
    2204.687, 2191.358, 2189.202, 2179.97, 2177.448, 2170.539, 2164.881, 
    2170.049, 2175.526, 2191.363, 2206.008, 2221.908, 2225.867, 2245.167, 
    2229.409, 2255.656, 2233.269, 2272.596, 2203.702, 2232.62, 2180.605, 
    2186.075, 2196.103, 2219.343, 2206.84, 2221.488, 2189.118, 2172.77, 
    2168.612, 2160.935, 2168.788, 2168.146, 2175.752, 2173.297, 2191.896, 
    2181.832, 2210.733, 2221.371, 2252.533, 2272.518, 2293.605, 2303.17, 
    2306.114, 2307.349,
  5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692,
  8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.706968, 4.725432, 4.721838, 4.73676, 4.728478, 4.738255, 4.710706, 
    4.726167, 4.716293, 4.708627, 4.765809, 4.737426, 4.795402, 4.777215, 
    4.822985, 4.79257, 4.829132, 4.822104, 4.843273, 4.837202, 4.864348, 
    4.846076, 4.878455, 4.85998, 4.862868, 4.845475, 4.743127, 4.76227, 
    4.741995, 4.744721, 4.743497, 4.72865, 4.72118, 4.705557, 4.708391, 
    4.719866, 4.745947, 4.737082, 4.759442, 4.758936, 4.783911, 4.77264, 
    4.814744, 4.802752, 4.837455, 4.828713, 4.837045, 4.834517, 4.837078, 
    4.82426, 4.829749, 4.81848, 4.77475, 4.787575, 4.749391, 4.726532, 
    4.711384, 4.700656, 4.702172, 4.705062, 4.719933, 4.733942, 4.744636, 
    4.751799, 4.758863, 4.780295, 4.791659, 4.817172, 4.812559, 4.820374, 
    4.827844, 4.840405, 4.838336, 4.843875, 4.820166, 4.835916, 4.809934, 
    4.817031, 4.760792, 4.739472, 4.730435, 4.722529, 4.703338, 4.716586, 
    4.71136, 4.723797, 4.731711, 4.727796, 4.751995, 4.742577, 4.792333, 
    4.77086, 4.826972, 4.813506, 4.830203, 4.821678, 4.836292, 4.823138, 
    4.845937, 4.850912, 4.847512, 4.860577, 4.82241, 4.837046, 4.727686, 
    4.728325, 4.731299, 4.718233, 4.717434, 4.70548, 4.716115, 4.720649, 
    4.73217, 4.738995, 4.745488, 4.759785, 4.775787, 4.79822, 4.814378, 
    4.825229, 4.818573, 4.824449, 4.817881, 4.814804, 4.849048, 4.829801, 
    4.858696, 4.857094, 4.844007, 4.857275, 4.728773, 4.725099, 4.712361, 
    4.722328, 4.704179, 4.714333, 4.720179, 4.742775, 4.747748, 4.752365, 
    4.761489, 4.773216, 4.793836, 4.811822, 4.828278, 4.827071, 4.827496, 
    4.831178, 4.822062, 4.832675, 4.834458, 4.829798, 4.85688, 4.849133, 
    4.85706, 4.852015, 4.726293, 4.732476, 4.729135, 4.73542, 4.730992, 
    4.750706, 4.756627, 4.784397, 4.772985, 4.791153, 4.774828, 4.777719, 
    4.79175, 4.775709, 4.810831, 4.787004, 4.831321, 4.807465, 4.832819, 
    4.828207, 4.835843, 4.842689, 4.851309, 4.867243, 4.86355, 4.876893, 
    4.741704, 4.749743, 4.749033, 4.757454, 4.763689, 4.777218, 4.798972, 
    4.790783, 4.805821, 4.808845, 4.786, 4.800019, 4.755127, 4.762362, 
    4.758053, 4.742338, 4.792671, 4.766798, 4.814646, 4.800575, 4.841713, 
    4.821228, 4.861518, 4.878811, 4.895114, 4.914218, 4.754133, 4.748666, 
    4.758456, 4.772025, 4.784634, 4.801433, 4.803153, 4.806306, 4.814476, 
    4.821353, 4.807304, 4.823078, 4.764044, 4.794921, 4.746602, 4.761119, 
    4.771224, 4.766788, 4.789848, 4.795294, 4.817466, 4.805995, 4.87454, 
    4.844138, 4.928791, 4.905042, 4.746758, 4.754113, 4.779775, 4.767553, 
    4.802555, 4.811197, 4.818228, 4.827229, 4.8282, 4.833538, 4.824792, 
    4.833192, 4.801469, 4.815629, 4.776835, 4.786259, 4.781922, 4.777168, 
    4.79185, 4.807525, 4.807858, 4.812892, 4.827101, 4.802697, 4.878477, 
    4.831592, 4.762143, 4.776351, 4.77838, 4.772872, 4.81033, 4.796736, 
    4.833407, 4.823478, 4.839753, 4.831662, 4.830472, 4.820094, 4.81364, 
    4.797359, 4.784139, 4.773671, 4.776103, 4.787606, 4.808485, 4.828289, 
    4.823946, 4.838515, 4.800012, 4.816134, 4.809899, 4.826167, 4.790566, 
    4.820878, 4.782839, 4.786166, 4.796466, 4.81723, 4.821828, 4.826746, 
    4.82371, 4.809015, 4.80661, 4.796216, 4.793349, 4.785441, 4.778902, 
    4.784877, 4.791158, 4.809021, 4.825156, 4.842787, 4.847107, 4.867776, 
    4.850949, 4.87874, 4.855111, 4.896057, 4.822635, 4.854413, 4.796935, 
    4.803105, 4.814281, 4.839973, 4.82609, 4.842328, 4.806515, 4.788005, 
    4.78322, 4.774307, 4.783424, 4.782682, 4.791417, 4.788609, 4.809614, 
    4.798324, 4.830443, 4.842199, 4.875494, 4.895977, 4.91688, 4.926127, 
    4.928943, 4.930121,
  6.780727, 6.803227, 6.798849, 6.817023, 6.806937, 6.818844, 6.785284, 
    6.804122, 6.792092, 6.78275, 6.852379, 6.817835, 6.88836, 6.866251, 
    6.921864, 6.884918, 6.929327, 6.920794, 6.946488, 6.939122, 6.97205, 
    6.94989, 6.98915, 6.966753, 6.970255, 6.94916, 6.824776, 6.848073, 
    6.823398, 6.826716, 6.825226, 6.807147, 6.798048, 6.779008, 6.782462, 
    6.796446, 6.828209, 6.817415, 6.844632, 6.844017, 6.874393, 6.860687, 
    6.911857, 6.897291, 6.939429, 6.928818, 6.938931, 6.935863, 6.938971, 
    6.923412, 6.930076, 6.916394, 6.863253, 6.878847, 6.832401, 6.804567, 
    6.78611, 6.773033, 6.774881, 6.778405, 6.796528, 6.813591, 6.826613, 
    6.835331, 6.843928, 6.869996, 6.883811, 6.914806, 6.909204, 6.918694, 
    6.927763, 6.943008, 6.940497, 6.947219, 6.918441, 6.93756, 6.906015, 
    6.914635, 6.846275, 6.820326, 6.809321, 6.799691, 6.776302, 6.792449, 
    6.786081, 6.801235, 6.810875, 6.806106, 6.83557, 6.824107, 6.88463, 
    6.858522, 6.926705, 6.910353, 6.930627, 6.920277, 6.938017, 6.92205, 
    6.949721, 6.955755, 6.951632, 6.967477, 6.921166, 6.938931, 6.805973, 
    6.806751, 6.810374, 6.794456, 6.793482, 6.778913, 6.791875, 6.7974, 
    6.811434, 6.819745, 6.82765, 6.845049, 6.864514, 6.891784, 6.911413, 
    6.924589, 6.916507, 6.923642, 6.915667, 6.91193, 6.953495, 6.930139, 
    6.965197, 6.963254, 6.947379, 6.963473, 6.807297, 6.802822, 6.787302, 
    6.799446, 6.777328, 6.789704, 6.796827, 6.824348, 6.830401, 6.83602, 
    6.847123, 6.861388, 6.886456, 6.908309, 6.92829, 6.926825, 6.927341, 
    6.93181, 6.920744, 6.933628, 6.935792, 6.930135, 6.962994, 6.953598, 
    6.963213, 6.957094, 6.804276, 6.811807, 6.807737, 6.815392, 6.809999, 
    6.834002, 6.841208, 6.874983, 6.861108, 6.883196, 6.863349, 6.866864, 
    6.883921, 6.86442, 6.907104, 6.878152, 6.931984, 6.903016, 6.933802, 
    6.928204, 6.937472, 6.94578, 6.956238, 6.97556, 6.971082, 6.987257, 
    6.823043, 6.832829, 6.831965, 6.842214, 6.849799, 6.866255, 6.892697, 
    6.882746, 6.90102, 6.904692, 6.876932, 6.89397, 6.839382, 6.848186, 
    6.842942, 6.823816, 6.885041, 6.853581, 6.911738, 6.894646, 6.944595, 
    6.919731, 6.968619, 6.989582, 7.009335, 7.032467, 6.838172, 6.831519, 
    6.843433, 6.85994, 6.875271, 6.895688, 6.897778, 6.901608, 6.911532, 
    6.919883, 6.902821, 6.921978, 6.850232, 6.887775, 6.829006, 6.846673, 
    6.858965, 6.85357, 6.881609, 6.888228, 6.915163, 6.90123, 6.984406, 
    6.947537, 7.050103, 7.021358, 6.829195, 6.838148, 6.869363, 6.8545, 
    6.897051, 6.907549, 6.916089, 6.927016, 6.928195, 6.934675, 6.924059, 
    6.934255, 6.895731, 6.912931, 6.865789, 6.877247, 6.871974, 6.866194, 
    6.884042, 6.90309, 6.903494, 6.909609, 6.926861, 6.897224, 6.989177, 
    6.932312, 6.847919, 6.865201, 6.867668, 6.86097, 6.906497, 6.889981, 
    6.934516, 6.922463, 6.942217, 6.932397, 6.930954, 6.918354, 6.910516, 
    6.890738, 6.874669, 6.861941, 6.864899, 6.878885, 6.904255, 6.928303, 
    6.923032, 6.940715, 6.893961, 6.913545, 6.905973, 6.925727, 6.882483, 
    6.919306, 6.87309, 6.877134, 6.889653, 6.914876, 6.92046, 6.92643, 
    6.922745, 6.904899, 6.901977, 6.889348, 6.885865, 6.876253, 6.868302, 
    6.875567, 6.883202, 6.904906, 6.9245, 6.945899, 6.95114, 6.976206, 
    6.955801, 6.989495, 6.960848, 7.010476, 6.921439, 6.960001, 6.890222, 
    6.89772, 6.911295, 6.942484, 6.925634, 6.945342, 6.901862, 6.879369, 
    6.873553, 6.862715, 6.873801, 6.872899, 6.883516, 6.880103, 6.905627, 
    6.89191, 6.930918, 6.945185, 6.985562, 7.01038, 7.035689, 7.04688, 
    7.050288, 7.051713,
  10.29747, 10.32977, 10.32348, 10.34957, 10.33509, 10.35218, 10.30401, 
    10.33105, 10.31378, 10.30037, 10.40032, 10.35073, 10.45198, 10.42024, 
    10.50008, 10.44704, 10.5108, 10.49854, 10.53544, 10.52486, 10.57214, 
    10.54032, 10.5967, 10.56453, 10.56956, 10.53927, 10.3607, 10.39414, 
    10.35872, 10.36348, 10.36135, 10.33539, 10.32233, 10.295, 10.29996, 
    10.32003, 10.36563, 10.35013, 10.3892, 10.38832, 10.43193, 10.41225, 
    10.48571, 10.4648, 10.5253, 10.51007, 10.52458, 10.52018, 10.52464, 
    10.5023, 10.51187, 10.49223, 10.41593, 10.43832, 10.37164, 10.33169, 
    10.3052, 10.28643, 10.28908, 10.29414, 10.32015, 10.34464, 10.36334, 
    10.37585, 10.38819, 10.42561, 10.44545, 10.48995, 10.4819, 10.49553, 
    10.50855, 10.53044, 10.52683, 10.53648, 10.49517, 10.52262, 10.47732, 
    10.4897, 10.39156, 10.35431, 10.33851, 10.32469, 10.29112, 10.31429, 
    10.30515, 10.32691, 10.34074, 10.3339, 10.37619, 10.35974, 10.44662, 
    10.40914, 10.50703, 10.48355, 10.51266, 10.4978, 10.52327, 10.50035, 
    10.54008, 10.54874, 10.54282, 10.56557, 10.49908, 10.52459, 10.33371, 
    10.33482, 10.34002, 10.31718, 10.31578, 10.29487, 10.31347, 10.3214, 
    10.34155, 10.35348, 10.36482, 10.3898, 10.41774, 10.45689, 10.48507, 
    10.50399, 10.49239, 10.50263, 10.49118, 10.48582, 10.5455, 10.51196, 
    10.5623, 10.55951, 10.53671, 10.55982, 10.33561, 10.32918, 10.30691, 
    10.32434, 10.29259, 10.31035, 10.32058, 10.36008, 10.36877, 10.37684, 
    10.39278, 10.41326, 10.44924, 10.48062, 10.50931, 10.5072, 10.50794, 
    10.51436, 10.49847, 10.51697, 10.52008, 10.51196, 10.55914, 10.54564, 
    10.55945, 10.55066, 10.33127, 10.34208, 10.33624, 10.34723, 10.33949, 
    10.37394, 10.38429, 10.43277, 10.41285, 10.44456, 10.41607, 10.42112, 
    10.44561, 10.41761, 10.47889, 10.43732, 10.51461, 10.47302, 10.51722, 
    10.50918, 10.52249, 10.53442, 10.54943, 10.57718, 10.57075, 10.59398, 
    10.35821, 10.37226, 10.37102, 10.38573, 10.39662, 10.42024, 10.45821, 
    10.44392, 10.47015, 10.47542, 10.43557, 10.46003, 10.38167, 10.3943, 
    10.38678, 10.35932, 10.44721, 10.40205, 10.48554, 10.461, 10.53272, 
    10.49702, 10.56721, 10.59731, 10.62568, 10.65891, 10.37993, 10.37038, 
    10.38748, 10.41118, 10.43319, 10.4625, 10.4655, 10.471, 10.48525, 
    10.49724, 10.47274, 10.50024, 10.39724, 10.45114, 10.36677, 10.39213, 
    10.40978, 10.40203, 10.44229, 10.45179, 10.49046, 10.47046, 10.58988, 
    10.53694, 10.68423, 10.64295, 10.36704, 10.37989, 10.42471, 10.40337, 
    10.46446, 10.47953, 10.49179, 10.50748, 10.50917, 10.51847, 10.50323, 
    10.51787, 10.46256, 10.48726, 10.41957, 10.43602, 10.42845, 10.42016, 
    10.44578, 10.47312, 10.47371, 10.48248, 10.50725, 10.4647, 10.59674, 
    10.51508, 10.39392, 10.41873, 10.42227, 10.41266, 10.47802, 10.4543, 
    10.51825, 10.50094, 10.5293, 10.5152, 10.51313, 10.49504, 10.48379, 
    10.45539, 10.43232, 10.41405, 10.4183, 10.43837, 10.4748, 10.50933, 
    10.50176, 10.52715, 10.46002, 10.48814, 10.47726, 10.50563, 10.44354, 
    10.49641, 10.43005, 10.43586, 10.45383, 10.49005, 10.49806, 10.50664, 
    10.50135, 10.47572, 10.47153, 10.4534, 10.4484, 10.4346, 10.42318, 
    10.43361, 10.44457, 10.47573, 10.50387, 10.53459, 10.54212, 10.57811, 
    10.54881, 10.59719, 10.55606, 10.62732, 10.49947, 10.55484, 10.45465, 
    10.46542, 10.48491, 10.52969, 10.50549, 10.53379, 10.47136, 10.43907, 
    10.43072, 10.41516, 10.43108, 10.42978, 10.44502, 10.44012, 10.47677, 
    10.45707, 10.51308, 10.53356, 10.59154, 10.62718, 10.66353, 10.67961, 
    10.6845, 10.68655,
  16.38583, 16.43753, 16.42747, 16.46924, 16.44606, 16.47342, 16.3963, 
    16.43958, 16.41194, 16.39048, 16.55055, 16.47111, 16.63338, 16.58248, 
    16.71057, 16.62545, 16.72777, 16.7081, 16.76734, 16.75035, 16.82631, 
    16.77518, 16.86578, 16.81409, 16.82217, 16.7735, 16.48706, 16.54065, 
    16.4839, 16.49153, 16.4881, 16.44654, 16.42562, 16.38188, 16.38981, 
    16.42194, 16.49496, 16.47014, 16.53273, 16.53132, 16.60122, 16.56967, 
    16.68751, 16.65395, 16.75106, 16.7266, 16.74991, 16.74284, 16.75, 
    16.71414, 16.7295, 16.69796, 16.57558, 16.61147, 16.5046, 16.44061, 
    16.3982, 16.36816, 16.3724, 16.3805, 16.42213, 16.46135, 16.49129, 
    16.51134, 16.53111, 16.5911, 16.6229, 16.6943, 16.68139, 16.70326, 
    16.72416, 16.75931, 16.75352, 16.76902, 16.70268, 16.74675, 16.67405, 
    16.69391, 16.53651, 16.47683, 16.45153, 16.4294, 16.37567, 16.41276, 
    16.39813, 16.43295, 16.45511, 16.44415, 16.51189, 16.48553, 16.62479, 
    16.56469, 16.72173, 16.68404, 16.73077, 16.70691, 16.7478, 16.711, 
    16.77479, 16.78871, 16.7792, 16.81576, 16.70896, 16.74991, 16.44384, 
    16.44563, 16.45395, 16.41737, 16.41513, 16.38166, 16.41144, 16.42414, 
    16.45639, 16.4755, 16.49367, 16.53369, 16.57848, 16.64127, 16.68648, 
    16.71685, 16.69822, 16.71466, 16.69629, 16.68767, 16.7835, 16.72964, 
    16.8105, 16.80601, 16.76939, 16.80652, 16.44688, 16.4366, 16.40093, 
    16.42884, 16.37802, 16.40645, 16.42282, 16.48608, 16.5, 16.51292, 
    16.53846, 16.57129, 16.62899, 16.67933, 16.72538, 16.722, 16.72319, 
    16.73349, 16.70799, 16.73768, 16.74267, 16.72963, 16.80541, 16.78374, 
    16.80592, 16.7918, 16.43994, 16.45725, 16.44789, 16.46549, 16.45309, 
    16.50828, 16.52485, 16.60258, 16.57064, 16.62149, 16.5758, 16.58389, 
    16.62316, 16.57827, 16.67656, 16.60987, 16.73389, 16.66714, 16.73808, 
    16.72518, 16.74655, 16.7657, 16.78983, 16.83441, 16.82408, 16.86141, 
    16.48308, 16.50558, 16.5036, 16.52717, 16.54462, 16.58249, 16.64337, 
    16.62045, 16.66254, 16.671, 16.60707, 16.6463, 16.52066, 16.54091, 
    16.52884, 16.48486, 16.62574, 16.55332, 16.68723, 16.64786, 16.76297, 
    16.70565, 16.81839, 16.86678, 16.91239, 16.96585, 16.51787, 16.50257, 
    16.52997, 16.56795, 16.60324, 16.65026, 16.65507, 16.66389, 16.68676, 
    16.706, 16.66669, 16.71083, 16.54562, 16.63203, 16.49679, 16.53743, 
    16.56571, 16.5533, 16.61783, 16.63308, 16.69512, 16.66302, 16.85483, 
    16.76976, 17.00662, 16.94017, 16.49723, 16.51782, 16.58964, 16.55544, 
    16.6534, 16.67758, 16.69726, 16.72244, 16.72516, 16.7401, 16.71563, 
    16.73913, 16.65036, 16.68998, 16.58142, 16.60779, 16.59565, 16.58235, 
    16.62344, 16.66731, 16.66824, 16.68233, 16.72208, 16.6538, 16.86584, 
    16.73465, 16.54029, 16.58006, 16.58574, 16.57032, 16.67516, 16.63711, 
    16.73973, 16.71195, 16.75749, 16.73485, 16.73152, 16.70248, 16.68442, 
    16.63886, 16.60186, 16.57256, 16.57937, 16.61156, 16.66999, 16.72541, 
    16.71326, 16.75402, 16.64628, 16.6914, 16.67395, 16.71947, 16.61985, 
    16.70467, 16.59822, 16.60753, 16.63636, 16.69446, 16.70733, 16.72109, 
    16.7126, 16.67147, 16.66474, 16.63565, 16.62763, 16.6055, 16.5872, 
    16.60392, 16.6215, 16.67149, 16.71664, 16.76598, 16.77807, 16.8359, 
    16.78882, 16.86658, 16.80046, 16.91503, 16.70959, 16.79851, 16.63767, 
    16.65494, 16.68621, 16.7581, 16.71926, 16.76469, 16.66448, 16.61268, 
    16.59929, 16.57434, 16.59986, 16.59778, 16.62222, 16.61437, 16.67315, 
    16.64155, 16.73144, 16.76433, 16.85749, 16.91481, 16.9733, 16.99917, 
    17.00705, 17.01035,
  26.07269, 26.16245, 26.14497, 26.21757, 26.17727, 26.22484, 26.09085, 
    26.16603, 26.11801, 26.08075, 26.35908, 26.22081, 26.50349, 26.41471, 
    26.63833, 26.48966, 26.66842, 26.63402, 26.73767, 26.70793, 26.841, 
    26.75141, 26.91025, 26.81957, 26.83374, 26.74846, 26.24856, 26.34182, 
    26.24305, 26.25632, 26.25037, 26.1781, 26.14177, 26.06583, 26.0796, 
    26.13538, 26.2623, 26.21913, 26.32804, 26.32557, 26.44738, 26.39239, 
    26.59802, 26.5394, 26.70917, 26.66637, 26.70716, 26.69478, 26.70732, 
    26.64458, 26.67144, 26.61629, 26.40268, 26.46527, 26.27907, 26.1678, 
    26.09415, 26.04202, 26.04939, 26.06343, 26.13571, 26.20385, 26.25591, 
    26.2908, 26.32522, 26.42974, 26.48521, 26.6099, 26.58734, 26.62556, 
    26.66211, 26.72362, 26.71348, 26.74062, 26.62454, 26.70163, 26.5745, 
    26.60921, 26.33462, 26.23077, 26.18679, 26.14833, 26.05505, 26.11943, 
    26.09403, 26.1545, 26.193, 26.17395, 26.29175, 26.24589, 26.4885, 
    26.38371, 26.65785, 26.59197, 26.67366, 26.63194, 26.70347, 26.63908, 
    26.75072, 26.7751, 26.75844, 26.8225, 26.63552, 26.70716, 26.17342, 
    26.17652, 26.19099, 26.12744, 26.12355, 26.06546, 26.11714, 26.13919, 
    26.19523, 26.22845, 26.26006, 26.32971, 26.40774, 26.51726, 26.59623, 
    26.64931, 26.61675, 26.6455, 26.61337, 26.59832, 26.76597, 26.67169, 
    26.81328, 26.80542, 26.74127, 26.8063, 26.1787, 26.16083, 26.0989, 
    26.14735, 26.05914, 26.10848, 26.1369, 26.24685, 26.27107, 26.29355, 
    26.33802, 26.3952, 26.49584, 26.58373, 26.66424, 26.65833, 26.66041, 
    26.67843, 26.63382, 26.68576, 26.6945, 26.67168, 26.80437, 26.76639, 
    26.80525, 26.78051, 26.16664, 26.19672, 26.18046, 26.21105, 26.1895, 
    26.28547, 26.31432, 26.44976, 26.39408, 26.48274, 26.40306, 26.41717, 
    26.48565, 26.40736, 26.57889, 26.46248, 26.67913, 26.56243, 26.68647, 
    26.66389, 26.70127, 26.73481, 26.77705, 26.8552, 26.83708, 26.90257, 
    26.24163, 26.28078, 26.27733, 26.31835, 26.34874, 26.41472, 26.52093, 
    26.48094, 26.5544, 26.56918, 26.45758, 26.52604, 26.30701, 26.34228, 
    26.32127, 26.24472, 26.49015, 26.3639, 26.59754, 26.52876, 26.73003, 
    26.62974, 26.82712, 26.91199, 26.99211, 27.08611, 26.30217, 26.27554, 
    26.32323, 26.38939, 26.45091, 26.53296, 26.54136, 26.55677, 26.59671, 
    26.63035, 26.56165, 26.63879, 26.35047, 26.50114, 26.26548, 26.33622, 
    26.38548, 26.36385, 26.47637, 26.50296, 26.61133, 26.55525, 26.89102, 
    26.74191, 27.15789, 27.04094, 26.26624, 26.30207, 26.4272, 26.36758, 
    26.53844, 26.58068, 26.61506, 26.6591, 26.66385, 26.68999, 26.64718, 
    26.68829, 26.53313, 26.60235, 26.41286, 26.45885, 26.43768, 26.41448, 
    26.48614, 26.56273, 26.56436, 26.58897, 26.65847, 26.53913, 26.91035, 
    26.68046, 26.34121, 26.41049, 26.42039, 26.39352, 26.57644, 26.51001, 
    26.68935, 26.64075, 26.72043, 26.6808, 26.67498, 26.62419, 26.59262, 
    26.51305, 26.44849, 26.39742, 26.40928, 26.46542, 26.56742, 26.66429, 
    26.64304, 26.71436, 26.52601, 26.60482, 26.57433, 26.6539, 26.47988, 
    26.62802, 26.44215, 26.45839, 26.50869, 26.61018, 26.63268, 26.65674, 
    26.64189, 26.57001, 26.55825, 26.50746, 26.49347, 26.45485, 26.42294, 
    26.4521, 26.48276, 26.57004, 26.64896, 26.73529, 26.75646, 26.85782, 
    26.77529, 26.91164, 26.79569, 26.99674, 26.63662, 26.79227, 26.51098, 
    26.54113, 26.59576, 26.7215, 26.65353, 26.73304, 26.55779, 26.46737, 
    26.44401, 26.40052, 26.44501, 26.44139, 26.48403, 26.47032, 26.57294, 
    26.51776, 26.67484, 26.73241, 26.89571, 26.99636, 27.09921, 27.14476, 
    27.15864, 27.16445,
  44.59721, 44.76149, 44.72948, 44.86251, 44.78864, 44.87585, 44.63044, 
    44.76804, 44.68012, 44.61195, 45.12243, 44.86846, 45.3885, 45.22482, 
    45.63772, 45.36298, 45.69342, 45.62974, 45.8218, 45.76664, 46.01373, 
    45.84729, 46.1426, 45.97388, 46.00022, 45.84182, 44.91938, 45.09069, 
    44.90926, 44.93362, 44.92268, 44.79016, 44.72362, 44.58468, 44.60986, 
    44.71191, 44.94458, 44.86538, 45.06535, 45.06082, 45.28503, 45.18372, 
    45.56313, 45.4548, 45.76894, 45.68962, 45.76522, 45.74227, 45.76551, 
    45.64927, 45.69902, 45.59693, 45.20267, 45.318, 44.97538, 44.77129, 
    44.63646, 44.54117, 44.55462, 44.58029, 44.71251, 44.83736, 44.93286, 
    44.99692, 45.06017, 45.2525, 45.35477, 45.5851, 45.54338, 45.61407, 
    45.68174, 45.79573, 45.77694, 45.82727, 45.61219, 45.75496, 45.51965, 
    45.58382, 45.07745, 44.88673, 44.80608, 44.73563, 44.56497, 44.68272, 
    44.63625, 44.74692, 44.81746, 44.78255, 44.99867, 44.91446, 45.36085, 
    45.16774, 45.67384, 45.55194, 45.70314, 45.62588, 45.75838, 45.63911, 
    45.84602, 45.89128, 45.86034, 45.97933, 45.63251, 45.76522, 44.78157, 
    44.78727, 44.81379, 44.69738, 44.69027, 44.584, 44.67853, 44.71889, 
    44.82156, 44.88246, 44.94047, 45.06842, 45.21199, 45.41391, 45.55983, 
    45.65805, 45.59777, 45.65098, 45.59151, 45.56368, 45.87432, 45.69949, 
    45.96218, 45.94759, 45.82847, 45.94923, 44.79126, 44.75852, 44.64515, 
    44.73384, 44.57244, 44.66268, 44.7147, 44.91623, 44.96068, 45.00198, 
    45.08369, 45.1889, 45.37438, 45.53671, 45.68568, 45.67474, 45.67859, 
    45.71198, 45.62937, 45.72556, 45.74174, 45.69946, 45.94563, 45.87509, 
    45.94727, 45.90132, 44.76916, 44.82429, 44.79449, 44.85056, 44.81105, 
    44.98714, 45.04014, 45.2894, 45.18683, 45.35022, 45.20338, 45.22935, 
    45.35559, 45.2113, 45.52775, 45.31285, 45.71327, 45.49734, 45.72686, 
    45.68504, 45.75431, 45.81649, 45.8949, 46.04014, 46.00644, 46.12831, 
    44.90666, 44.97852, 44.97218, 45.04755, 45.10341, 45.22485, 45.42069, 
    45.34689, 45.4825, 45.50981, 45.30382, 45.43013, 45.02671, 45.09152, 
    45.05291, 44.91233, 45.36389, 45.13129, 45.56224, 45.43515, 45.80762, 
    45.6218, 45.98791, 46.14586, 46.29525, 46.47086, 45.0178, 44.96889, 
    45.05652, 45.1782, 45.29153, 45.44289, 45.45842, 45.48688, 45.56071, 
    45.62294, 45.49589, 45.63856, 45.1066, 45.38417, 44.95043, 45.08038, 
    45.17101, 45.13121, 45.33846, 45.38753, 45.58776, 45.48407, 46.10681, 
    45.82966, 46.60526, 46.38643, 44.95182, 45.01763, 45.24783, 45.13807, 
    45.45302, 45.53107, 45.59466, 45.67617, 45.68497, 45.73338, 45.65409, 
    45.73024, 45.44321, 45.57113, 45.22141, 45.30616, 45.26714, 45.2244, 
    45.35649, 45.49789, 45.5009, 45.54639, 45.675, 45.4543, 46.14281, 
    45.71572, 45.08956, 45.21706, 45.2353, 45.18581, 45.52323, 45.40053, 
    45.7322, 45.64219, 45.78981, 45.71637, 45.70557, 45.61154, 45.55315, 
    45.40615, 45.28707, 45.19298, 45.21483, 45.31828, 45.50656, 45.68578, 
    45.64643, 45.77857, 45.43007, 45.57571, 45.51934, 45.66654, 45.34493, 
    45.61863, 45.27539, 45.30532, 45.3981, 45.58562, 45.62725, 45.67179, 
    45.64429, 45.51135, 45.48962, 45.39583, 45.37, 45.2988, 45.23999, 
    45.29372, 45.35026, 45.5114, 45.65739, 45.81738, 45.85666, 46.04501, 
    45.89162, 46.14521, 45.92951, 46.30389, 45.63454, 45.92315, 45.40232, 
    45.45798, 45.55895, 45.79181, 45.66585, 45.81321, 45.48877, 45.32187, 
    45.27882, 45.1987, 45.28065, 45.27398, 45.35259, 45.3273, 45.51676, 
    45.41484, 45.70531, 45.81203, 46.11553, 46.30317, 46.49539, 46.58067, 
    46.60667, 46.61755,
  75.10475, 75.4586, 75.38952, 75.67706, 75.51723, 75.70596, 75.17618, 
    75.47274, 75.28311, 75.13644, 76.24215, 75.68993, 76.82531, 76.466, 
    77.37594, 76.76917, 77.49962, 77.35824, 77.78548, 77.66252, 78.21509, 
    77.84238, 78.5051, 78.12568, 78.18476, 77.83015, 75.80031, 76.17292, 
    75.77837, 75.83121, 75.80749, 75.52055, 75.37688, 75.07784, 75.13192, 
    75.35164, 75.85501, 75.68327, 76.11768, 76.10781, 76.59796, 76.37608, 
    77.21069, 76.97137, 77.66764, 77.49117, 77.65934, 77.60825, 77.66, 
    77.40157, 77.51205, 77.28553, 76.41753, 76.67033, 75.92191, 75.47976, 
    75.18914, 74.98443, 75.01329, 75.0684, 75.35294, 75.6226, 75.82957, 
    75.96873, 76.10639, 76.52665, 76.75113, 77.25932, 77.167, 77.32352, 
    77.47367, 77.72734, 77.68545, 77.79769, 77.31935, 77.63651, 77.11454, 
    77.2565, 76.14404, 75.72952, 75.55495, 75.40279, 75.03551, 75.28873, 
    75.18868, 75.42715, 75.57957, 75.5041, 75.97253, 75.78966, 76.76448, 
    76.34114, 77.45612, 77.18593, 77.5212, 77.34969, 77.64411, 77.37902, 
    77.83955, 77.94069, 77.87154, 78.13789, 77.3644, 77.65935, 75.50199, 
    75.51428, 75.57162, 75.3203, 75.30499, 75.07635, 75.2797, 75.36668, 
    75.58841, 75.72028, 75.84609, 76.12437, 76.43792, 76.88126, 77.20338, 
    77.42105, 77.2874, 77.40536, 77.27353, 77.2119, 77.90276, 77.51309, 
    78.09946, 78.06673, 77.80037, 78.07042, 75.52292, 75.4522, 75.20783, 
    75.39893, 75.05155, 75.24557, 75.35764, 75.7935, 75.88998, 75.97973, 
    76.15766, 76.38741, 76.79425, 77.15226, 77.48242, 77.45811, 77.46667, 
    77.54086, 77.35742, 77.57106, 77.60706, 77.51303, 78.06236, 77.9045, 
    78.06604, 77.96315, 75.47517, 75.59432, 75.52989, 75.65117, 75.56569, 
    75.94746, 76.06277, 76.60755, 76.38287, 76.74112, 76.41908, 76.47593, 
    76.75292, 76.43639, 77.13245, 76.65903, 77.54374, 77.06526, 77.57395, 
    77.48099, 77.63504, 77.77364, 77.94878, 78.27444, 78.19874, 78.47289, 
    75.77273, 75.92873, 75.91495, 76.0789, 76.20067, 76.46607, 76.89619, 
    76.7338, 77.03249, 77.09279, 76.63921, 76.917, 76.03353, 76.17474, 
    76.09058, 75.78503, 76.77118, 76.26151, 77.20873, 76.92806, 77.75384, 
    77.34065, 78.15714, 78.51244, 78.85021, 79.24949, 76.01415, 75.90781, 
    76.09844, 76.36401, 76.61223, 76.94511, 76.97935, 77.04215, 77.20534, 
    77.34318, 77.06206, 77.37782, 76.20762, 76.81577, 75.86771, 76.15044, 
    76.34829, 76.26133, 76.71528, 76.82317, 77.26521, 77.03596, 78.42442, 
    77.80302, 79.55668, 79.05723, 75.87074, 76.01378, 76.5164, 76.27632, 
    76.96745, 77.13977, 77.28049, 77.46128, 77.48083, 77.58848, 77.41228, 
    77.58149, 76.94583, 77.2284, 76.45854, 76.64433, 76.55872, 76.46509, 
    76.75491, 77.06647, 77.07312, 77.17367, 77.4587, 76.97028, 78.50556, 
    77.54919, 76.17045, 76.44902, 76.48895, 76.38065, 77.12246, 76.85178, 
    77.58585, 77.38586, 77.71414, 77.55061, 77.52663, 77.31789, 77.18861, 
    76.86416, 76.60245, 76.39633, 76.44415, 76.67094, 77.08562, 77.48263, 
    77.39526, 77.68908, 76.91685, 77.23853, 77.11385, 77.43991, 76.7295, 
    77.33363, 76.57681, 76.64249, 76.84644, 77.26048, 77.35272, 77.45156, 
    77.39053, 77.0962, 77.04821, 76.84145, 76.78461, 76.62817, 76.49922, 
    76.61703, 76.7412, 77.09631, 77.41959, 77.77562, 77.8633, 78.28538, 
    77.94145, 78.51097, 78.02625, 78.86981, 77.3689, 78.01201, 76.85574, 
    76.97839, 77.20145, 77.7186, 77.43837, 77.7663, 77.04633, 76.67882, 
    76.58434, 76.40883, 76.58836, 76.57372, 76.74633, 76.69076, 77.10816, 
    76.88331, 77.52603, 77.76369, 78.44407, 78.86816, 79.30544, 79.50036, 
    79.55991, 79.58485,
  138.2295, 139.2781, 139.0721, 139.9332, 139.4533, 140.0204, 138.4399, 
    139.3203, 138.7561, 138.3228, 141.6568, 139.972, 143.4813, 142.3514, 
    145.2499, 143.3035, 145.6535, 145.1923, 146.5958, 146.1889, 148.0374, 
    146.785, 149.0286, 147.7348, 147.9347, 146.7443, 140.3055, 141.4433, 
    140.2391, 140.3992, 140.3273, 139.4632, 139.0345, 138.1504, 138.3095, 
    138.9595, 140.4714, 139.952, 141.2735, 141.2432, 142.7643, 142.0716, 
    144.7143, 143.946, 146.2058, 145.6259, 146.1784, 146.0101, 146.1806, 
    145.3333, 145.6942, 144.9563, 142.2004, 142.9917, 140.6748, 139.3413, 
    138.4782, 137.8764, 137.961, 138.1226, 138.9633, 139.7693, 140.3942, 
    140.8175, 141.2388, 142.5409, 143.2465, 144.8714, 144.5734, 145.0795, 
    145.5686, 146.4031, 146.2646, 146.6364, 145.066, 146.1031, 144.4046, 
    144.8623, 141.3545, 140.0914, 139.5663, 139.1116, 138.0261, 138.7728, 
    138.4768, 139.1842, 139.6401, 139.414, 140.8291, 140.2733, 143.2887, 
    141.9631, 145.5113, 144.6344, 145.7242, 145.1645, 146.1282, 145.2599, 
    146.7756, 147.1131, 146.8822, 147.7761, 145.2123, 146.1784, 139.4077, 
    139.4445, 139.6163, 138.8664, 138.821, 138.146, 138.746, 139.0042, 
    139.6666, 140.0636, 140.4444, 141.294, 142.2639, 143.6589, 144.6907, 
    145.3968, 144.9624, 145.3457, 144.9174, 144.7182, 146.9863, 145.6976, 
    147.6463, 147.5361, 146.6453, 147.5485, 139.4703, 139.259, 138.5334, 
    139.1001, 138.0732, 138.645, 138.9773, 140.2849, 140.5777, 140.8511, 
    141.3963, 142.1067, 143.3829, 144.5259, 145.5972, 145.5178, 145.5457, 
    145.7886, 145.1896, 145.8878, 146.0062, 145.6974, 147.5213, 146.9921, 
    147.5338, 147.1883, 139.3275, 139.6844, 139.4912, 139.8553, 139.5985, 
    140.7527, 141.105, 142.7944, 142.0927, 143.2149, 142.2053, 142.3824, 
    143.2522, 142.2592, 144.4621, 142.9561, 145.7981, 144.2464, 145.8973, 
    145.5925, 146.0983, 146.5565, 147.1402, 148.2391, 147.982, 148.9178, 
    140.2221, 140.6956, 140.6536, 141.1545, 141.5288, 142.3517, 143.7064, 
    143.1918, 144.1414, 144.3347, 142.8938, 143.7727, 141.0155, 141.4489, 
    141.1903, 140.2593, 143.3099, 141.7166, 144.7079, 143.8079, 146.4909, 
    145.1351, 147.8412, 149.0539, 150.2278, 151.6432, 140.9563, 140.6319, 
    141.2144, 142.0341, 142.8091, 143.8622, 143.9715, 144.1723, 144.697, 
    145.1433, 144.2361, 145.256, 141.5502, 143.4511, 140.51, 141.3741, 
    141.9853, 141.716, 143.1333, 143.4745, 144.8905, 144.1525, 148.7514, 
    146.6541, 152.7535, 150.9578, 140.5192, 140.9551, 142.5088, 141.7623, 
    143.9335, 144.4857, 144.94, 145.5281, 145.5921, 145.945, 145.3682, 
    145.922, 143.8645, 144.7715, 142.3282, 142.9099, 142.6413, 142.3486, 
    143.2585, 144.2503, 144.2716, 144.5948, 145.5197, 143.9425, 149.0302, 
    145.816, 141.4357, 142.2985, 142.4231, 142.0857, 144.43, 143.5653, 
    145.9364, 145.2821, 146.3595, 145.8206, 145.742, 145.0612, 144.643, 
    143.6046, 142.7783, 142.1345, 142.2833, 142.9936, 144.3117, 145.5979, 
    145.3128, 146.2766, 143.7722, 144.8042, 144.4023, 145.4583, 143.1782, 
    145.1123, 142.6979, 142.9041, 143.5483, 144.8752, 145.1743, 145.4964, 
    145.2973, 144.3456, 144.1917, 143.5325, 143.3524, 142.8591, 142.4551, 
    142.8241, 143.2152, 144.346, 145.392, 146.5631, 146.8547, 148.2763, 
    147.1156, 149.0488, 147.3999, 150.2966, 145.227, 147.3521, 143.5779, 
    143.9684, 144.6844, 146.3742, 145.4533, 146.5322, 144.1857, 143.0184, 
    142.7215, 142.1734, 142.7341, 142.6882, 143.2314, 143.056, 144.3841, 
    143.6655, 145.74, 146.5235, 148.8188, 150.2908, 151.844, 152.5485, 
    152.7653, 152.8563,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.01747908, -0.01720448, -0.0172575, -0.01703868, -0.0171597, -0.01701695, 
    -0.01742304, -0.01719367, -0.01733972, -0.01745418, -0.01662251, 
    -0.01702899, -0.0162115, -0.01646258, -0.01583977, -0.01625028, 
    -0.01575837, -0.01585148, -0.01557311, -0.01565231, -0.01530201, 
    -0.0155367, -0.01512384, -0.01535772, -0.01532086, -0.01554451, 
    -0.01694636, -0.01667253, -0.01696273, -0.01692335, -0.01694101, 
    -0.01715719, -0.01726723, -0.01750028, -0.01745773, -0.01728669, 
    -0.01690567, -0.017034, -0.01671263, -0.01671982, -0.01636957, 
    -0.0165265, -0.01594971, -0.01611139, -0.015649, -0.0157639, -0.01565437, 
    -0.0156875, -0.01565394, -0.01582284, -0.01575023, -0.01589975, 
    -0.01649698, -0.01631896, -0.01685614, -0.0171883, -0.01741291, 
    -0.01757419, -0.01755129, -0.01750772, -0.0172857, -0.01707975, 
    -0.01692457, -0.01682162, -0.01672085, -0.01641972, -0.01626278, 
    -0.01591722, -0.01597901, -0.0158745, -0.01577539, -0.01561047, 
    -0.01563749, -0.01556528, -0.01587727, -0.01566916, -0.01601432, 
    -0.01591909, -0.01669347, -0.01699928, -0.01713101, -0.0172473, 
    -0.01753371, -0.01733537, -0.01741326, -0.01722858, -0.01711233, 
    -0.01716972, -0.01681882, -0.0169543, -0.01625353, -0.01655145, 
    -0.01578691, -0.01596631, -0.01574424, -0.01585714, -0.01566423, 
    -0.01583773, -0.01553851, -0.01547416, -0.0155181, -0.01535009, 
    -0.01584741, -0.01565436, -0.01717133, -0.01716195, -0.01711835, 
    -0.01731091, -0.01732277, -0.01750145, -0.01734237, -0.0172751, 
    -0.01710562, -0.01700621, -0.01691229, -0.01670776, -0.01648249, 
    -0.01617303, -0.01595461, -0.01580999, -0.01589851, -0.01582033, 
    -0.01590775, -0.0159489, -0.01549823, -0.01574955, -0.01537413, 
    -0.01539465, -0.01556356, -0.01539234, -0.01715538, -0.01720938, 
    -0.01739831, -0.01725027, -0.01752103, -0.01736889, -0.01728206, 
    -0.01695144, -0.01687974, -0.01681353, -0.01668359, -0.01651842, 
    -0.01623294, -0.01598892, -0.01576965, -0.0157856, -0.01577998, 
    -0.0157314, -0.01585202, -0.0157117, -0.01568827, -0.01574959, 
    -0.0153974, -0.01549713, -0.01539509, -0.01545994, -0.01719181, 
    -0.01710114, -0.01715007, -0.01705818, -0.01712285, -0.01683728, 
    -0.01675267, -0.01636285, -0.01652165, -0.01626972, -0.01649588, 
    -0.01645555, -0.01626153, -0.01648358, -0.01600225, -0.01632684, 
    -0.01572952, -0.01604761, -0.01570981, -0.01577059, -0.01567011, 
    -0.01558071, -0.01546903, -0.01526524, -0.01531217, -0.01514344, 
    -0.01696694, -0.01685109, -0.01686128, -0.01674089, -0.01665245, 
    -0.01646253, -0.01616278, -0.01627481, -0.01606981, -0.01602899, 
    -0.01634069, -0.01614853, -0.01677405, -0.01667122, -0.01673238, 
    -0.01695776, -0.01624889, -0.01660857, -0.01595102, -0.01614096, 
    -0.01559342, -0.01586313, -0.01533807, -0.01511937, -0.01491673, 
    -0.01468358, -0.01678825, -0.01686655, -0.01672664, -0.01653511, 
    -0.01635957, -0.0161293, -0.01610595, -0.01606327, -0.01595329, 
    -0.01586146, -0.01604978, -0.01583853, -0.01664743, -0.01621808, 
    -0.01689624, -0.01668883, -0.01654634, -0.0166087, -0.01628767, 
    -0.01621298, -0.01591329, -0.01606746, -0.01517302, -0.01556187, 
    -0.01450878, -0.014795, -0.016894, -0.01678853, -0.01642695, -0.01659792, 
    -0.01611406, -0.01599732, -0.01590311, -0.01578352, -0.01577068, 
    -0.01570036, -0.01581578, -0.01570491, -0.01612881, -0.01593786, 
    -0.01646787, -0.01633712, -0.01639713, -0.01646323, -0.01626017, 
    -0.01604679, -0.01604229, -0.01597453, -0.01578521, -0.01611214, 
    -0.01512355, -0.01572595, -0.01667432, -0.01647461, -0.01644634, 
    -0.01652324, -0.01600898, -0.01619327, -0.01570207, -0.01583321, 
    -0.01561897, -0.01572503, -0.0157407, -0.01587823, -0.01596451, 
    -0.01618477, -0.01636643, -0.01651207, -0.01647808, -0.01631853, 
    -0.01603384, -0.01576951, -0.015827, -0.01563514, -0.01614863, 
    -0.0159311, -0.01601478, -0.01579757, -0.01627779, -0.01586779, 
    -0.01638441, -0.0163384, -0.01619696, -0.01591644, -0.01585514, 
    -0.01578991, -0.01583013, -0.01602669, -0.01605916, -0.01620039, 
    -0.0162396, -0.01634841, -0.01643908, -0.01635621, -0.01626966, 
    -0.01602662, -0.01581096, -0.01557943, -0.01552335, -0.01525847, 
    -0.01547368, -0.01512027, -0.0154201, -0.01490512, -0.01584442, 
    -0.01542908, -0.01619056, -0.0161066, -0.0159559, -0.0156161, 
    -0.01579859, -0.01558541, -0.01606044, -0.01631304, -0.01637913, 
    -0.01650317, -0.01637631, -0.01638659, -0.01626611, -0.01630472, 
    -0.01601862, -0.01617162, -0.01574109, -0.01558709, -0.01516102, 
    -0.0149061, -0.01465146, -0.01454054, -0.01450696, -0.01449295,
  -0.02241801, -0.02206922, -0.02213657, -0.0218586, -0.02201234, 
    -0.02183099, -0.02234684, -0.02205548, -0.02224101, -0.02238639, 
    -0.02132986, -0.02184629, -0.02080759, -0.02112665, -0.02033513, 
    -0.02085687, -0.02023166, -0.02035001, -0.01999616, -0.02009684, 
    -0.01965149, -0.01994988, -0.01942494, -0.01972233, -0.01967546, 
    -0.0199598, -0.02174132, -0.02139342, -0.02176211, -0.02171208, 
    -0.02173452, -0.02200914, -0.02214893, -0.02244494, -0.02239089, 
    -0.02217365, -0.02168962, -0.02185265, -0.02144437, -0.0214535, 
    -0.02100846, -0.02120787, -0.02047487, -0.02068036, -0.02009263, 
    -0.0202387, -0.02009946, -0.02014157, -0.02009891, -0.02031361, 
    -0.02022131, -0.02041137, -0.02117036, -0.02094414, -0.0216267, 
    -0.02204866, -0.02233396, -0.02253882, -0.02250973, -0.02245439, 
    -0.02217238, -0.02191077, -0.02171364, -0.02158284, -0.02145481, 
    -0.02107218, -0.02087275, -0.02043357, -0.02051211, -0.02037928, 
    -0.02025329, -0.02004365, -0.020078, -0.01998621, -0.02038279, 
    -0.02011826, -0.02055698, -0.02043596, -0.02142002, -0.02180855, 
    -0.02197589, -0.0221236, -0.0224874, -0.02223547, -0.02233441, 
    -0.02209984, -0.02195216, -0.02202507, -0.02157928, -0.02175141, 
    -0.020861, -0.02123957, -0.02026794, -0.02049596, -0.02021371, 
    -0.02035721, -0.02011199, -0.02033254, -0.01995217, -0.01987037, 
    -0.01992623, -0.01971262, -0.02034484, -0.02009945, -0.02202711, 
    -0.0220152, -0.02195981, -0.0222044, -0.02221947, -0.02244642, 
    -0.02224437, -0.02215892, -0.02194364, -0.02181735, -0.02169803, 
    -0.02143819, -0.02115196, -0.02075869, -0.0204811, -0.02029728, 
    -0.02040979, -0.02031042, -0.02042153, -0.02047384, -0.01990097, 
    -0.02022045, -0.01974319, -0.01976928, -0.01998402, -0.01976633, 
    -0.02200684, -0.02207545, -0.02231542, -0.02212738, -0.02247129, 
    -0.02227806, -0.02216776, -0.02174777, -0.02165669, -0.02157256, 
    -0.02140748, -0.02119761, -0.02083483, -0.0205247, -0.020246, 
    -0.02026628, -0.02025913, -0.02019738, -0.0203507, -0.02017233, 
    -0.02014255, -0.0202205, -0.01977277, -0.01989957, -0.01976983, 
    -0.01985228, -0.02205312, -0.02193795, -0.0220001, -0.02188337, 
    -0.02196553, -0.02160273, -0.02149523, -0.02099992, -0.02120171, 
    -0.02088158, -0.02116896, -0.02111772, -0.02087117, -0.02115333, 
    -0.02054165, -0.02095416, -0.02019499, -0.0205993, -0.02016994, 
    -0.02024719, -0.02011947, -0.02000581, -0.01986385, -0.01960474, 
    -0.01966441, -0.01944987, -0.02176746, -0.02162028, -0.02163322, 
    -0.02148028, -0.02136791, -0.02112659, -0.02074567, -0.02088804, 
    -0.02062752, -0.02057564, -0.02097177, -0.02072755, -0.02152241, 
    -0.02139175, -0.02146946, -0.0217558, -0.0208551, -0.02131216, 
    -0.02047654, -0.02071794, -0.02002197, -0.02036482, -0.01969734, 
    -0.01941927, -0.01916157, -0.01886505, -0.02154044, -0.02163993, 
    -0.02146217, -0.02121881, -0.02099575, -0.02070312, -0.02067344, 
    -0.02061919, -0.02047943, -0.0203627, -0.02060205, -0.02033355, 
    -0.02136152, -0.02081595, -0.02167764, -0.02141413, -0.02123308, 
    -0.02131232, -0.02090438, -0.02080947, -0.02042858, -0.02062453, 
    -0.01948748, -0.01998187, -0.01864271, -0.01900676, -0.0216748, 
    -0.0215408, -0.02108137, -0.02129862, -0.02068376, -0.02053538, 
    -0.02041563, -0.02026363, -0.02024731, -0.02015792, -0.02030463, 
    -0.0201637, -0.0207025, -0.02045981, -0.02113337, -0.02096722, 
    -0.02104349, -0.02112747, -0.02086943, -0.02059826, -0.02059254, 
    -0.02050642, -0.02026578, -0.0206813, -0.01942458, -0.02019046, 
    -0.0213957, -0.02114194, -0.02110601, -0.02120373, -0.0205502, 
    -0.02078442, -0.0201601, -0.0203268, -0.02005446, -0.02018928, 
    -0.0202092, -0.02038402, -0.02049368, -0.02077361, -0.02100447, 
    -0.02118953, -0.02114634, -0.0209436, -0.0205818, -0.02024582, 
    -0.0203189, -0.02007501, -0.02072768, -0.02045121, -0.02055757, 
    -0.0202815, -0.02089183, -0.02037074, -0.02102732, -0.02096885, 
    -0.0207891, -0.02043258, -0.02035466, -0.02027176, -0.02032288, 
    -0.02057271, -0.02061398, -0.02079346, -0.0208433, -0.02098157, 
    -0.02109679, -0.02099148, -0.0208815, -0.02057262, -0.02029851, 
    -0.0200042, -0.0199329, -0.01959614, -0.01986975, -0.0194204, 
    -0.01980164, -0.01914681, -0.02034104, -0.01981305, -0.02078097, 
    -0.02067427, -0.02048274, -0.02005081, -0.02028278, -0.02001179, 
    -0.0206156, -0.02093663, -0.02102061, -0.02117822, -0.02101703, 
    -0.02103009, -0.02087699, -0.02092605, -0.02056245, -0.0207569, 
    -0.02020969, -0.02001393, -0.01947222, -0.01914805, -0.01882419, 
    -0.0186831, -0.01864039, -0.01862257,
  -0.02349876, -0.02313152, -0.02320243, -0.02290973, -0.02307162, 
    -0.02288065, -0.02342382, -0.02311705, -0.0233124, -0.02346547, 
    -0.02235287, -0.02289676, -0.0218027, -0.02213882, -0.02130489, 
    -0.02185462, -0.02119586, -0.02132058, -0.02094767, -0.02105378, 
    -0.0205844, -0.0208989, -0.02034558, -0.02065906, -0.02060966, 
    -0.02090935, -0.02278621, -0.02241981, -0.02280812, -0.02275543, 
    -0.02277906, -0.02306825, -0.02321545, -0.02352711, -0.02347021, 
    -0.02324147, -0.02273178, -0.02290346, -0.02247348, -0.02248309, 
    -0.02201432, -0.02222436, -0.02145214, -0.02166865, -0.02104934, 
    -0.02120327, -0.02105654, -0.02110092, -0.02105596, -0.02128221, 
    -0.02118495, -0.02138523, -0.02218486, -0.02194656, -0.0226655, 
    -0.02310987, -0.02341027, -0.02362594, -0.02359532, -0.02353706, 
    -0.02324014, -0.02296466, -0.02275707, -0.02261932, -0.02248448, 
    -0.02208144, -0.02187135, -0.02140862, -0.02149138, -0.02135141, 
    -0.02121866, -0.02099772, -0.02103392, -0.02093718, -0.02135511, 
    -0.02107636, -0.02153866, -0.02141114, -0.02244783, -0.02285702, 
    -0.02303324, -0.02318878, -0.02357181, -0.02330657, -0.02341074, 
    -0.02316375, -0.02300825, -0.02308502, -0.02261556, -0.02279685, 
    -0.02185897, -0.02225777, -0.02123409, -0.02147437, -0.02117694, 
    -0.02132816, -0.02106975, -0.02130216, -0.02090131, -0.02081509, 
    -0.02087397, -0.02064883, -0.02131512, -0.02105653, -0.02308717, 
    -0.02307463, -0.02301631, -0.02327386, -0.02328972, -0.02352867, 
    -0.02331594, -0.02322596, -0.02299928, -0.02286628, -0.02274063, 
    -0.02246696, -0.02216547, -0.02175118, -0.0214587, -0.02126501, 
    -0.02138356, -0.02127886, -0.02139594, -0.02145106, -0.02084735, 
    -0.02118404, -0.02068105, -0.02070855, -0.02093488, -0.02070545, 
    -0.02306583, -0.02313807, -0.02339074, -0.02319276, -0.02355485, 
    -0.02335141, -0.02323528, -0.02279301, -0.02269709, -0.02260849, 
    -0.02243462, -0.02221356, -0.0218314, -0.02150464, -0.02121096, 
    -0.02123234, -0.02122481, -0.02115974, -0.0213213, -0.02113334, 
    -0.02110196, -0.0211841, -0.02071223, -0.02084588, -0.02070913, 
    -0.02079603, -0.02311457, -0.02299328, -0.02305873, -0.02293582, 
    -0.02302233, -0.02264027, -0.02252705, -0.02200532, -0.02221788, 
    -0.02188064, -0.02218338, -0.02212941, -0.02186968, -0.02216692, 
    -0.0215225, -0.02195711, -0.02115721, -0.02158324, -0.02113081, 
    -0.02121223, -0.02107763, -0.02095785, -0.02080822, -0.02053511, 
    -0.02059801, -0.02037186, -0.02281375, -0.02265875, -0.02267238, 
    -0.02251129, -0.02239295, -0.02213875, -0.02173747, -0.02188745, 
    -0.02161298, -0.02155832, -0.02197566, -0.02171838, -0.02255567, 
    -0.02241805, -0.0224999, -0.02280147, -0.02185276, -0.02233422, 
    -0.0214539, -0.02170824, -0.02097488, -0.02133618, -0.02063273, 
    -0.0203396, -0.02006792, -0.01975526, -0.02257466, -0.02267944, 
    -0.02249223, -0.02223589, -0.02200093, -0.02169263, -0.02166137, 
    -0.02160421, -0.02145694, -0.02133394, -0.02158615, -0.02130323, 
    -0.02238622, -0.0218115, -0.02271916, -0.02244162, -0.02225093, 
    -0.02233439, -0.02190467, -0.02180468, -0.02140336, -0.02160983, 
    -0.0204115, -0.02093261, -0.0195208, -0.01990469, -0.02271616, 
    -0.02257504, -0.02209112, -0.02231997, -0.02167223, -0.0215159, 
    -0.02138972, -0.02122955, -0.02121236, -0.02111815, -0.02127276, 
    -0.02112424, -0.02169198, -0.02143627, -0.02214589, -0.02197087, 
    -0.02205121, -0.02213968, -0.02186785, -0.02158215, -0.02157612, 
    -0.02148538, -0.02123182, -0.02166965, -0.0203452, -0.02115244, 
    -0.02242221, -0.02215492, -0.02211707, -0.02222001, -0.02153151, 
    -0.02177829, -0.02112045, -0.02129611, -0.02100911, -0.0211512, 
    -0.02117219, -0.02135641, -0.02147196, -0.0217669, -0.0220101, 
    -0.02220505, -0.02215956, -0.02194599, -0.02156481, -0.02121078, 
    -0.02128779, -0.02103078, -0.02171851, -0.02142721, -0.02153928, 
    -0.02124837, -0.02189144, -0.02134242, -0.02203418, -0.02197259, 
    -0.02178322, -0.02140758, -0.02132547, -0.02123811, -0.02129198, 
    -0.02155523, -0.02159871, -0.02178781, -0.02184032, -0.02198599, 
    -0.02210736, -0.02199643, -0.02188056, -0.02155514, -0.0212663, 
    -0.02095614, -0.020881, -0.02052605, -0.02081445, -0.02034079, 
    -0.02074266, -0.02005236, -0.02131112, -0.02075468, -0.02177466, 
    -0.02166224, -0.02146043, -0.02100527, -0.02124973, -0.02096415, 
    -0.02160042, -0.02193864, -0.02202712, -0.02219314, -0.02202334, 
    -0.0220371, -0.02187581, -0.0219275, -0.02154442, -0.0217493, 
    -0.02117271, -0.0209664, -0.02039542, -0.02005367, -0.01971218, 
    -0.0195634, -0.01951836, -0.01949956,
  -0.02299424, -0.02262573, -0.02269689, -0.02240317, -0.02256563, -0.022374, 
    -0.02291904, -0.02261121, -0.02280723, -0.02296083, -0.02184436, 
    -0.02239016, -0.02129221, -0.02162954, -0.02079258, -0.02134432, 
    -0.02068315, -0.02080832, -0.02043403, -0.02054054, -0.02006939, 
    -0.02038507, -0.01982967, -0.02014433, -0.02009475, -0.02039557, 
    -0.02227923, -0.02191154, -0.02230121, -0.02224833, -0.02227205, 
    -0.02256224, -0.02270995, -0.02302268, -0.02296558, -0.02273607, 
    -0.0222246, -0.02239689, -0.02196539, -0.02197504, -0.02150459, 
    -0.02171539, -0.02094037, -0.02115767, -0.02053608, -0.02069058, 
    -0.02054331, -0.02058785, -0.02054273, -0.02076982, -0.0206722, 
    -0.02087321, -0.02167574, -0.02143659, -0.0221581, -0.02260401, 
    -0.02290544, -0.02312185, -0.02309112, -0.02303267, -0.02273473, 
    -0.0224583, -0.02224998, -0.02211175, -0.02197643, -0.02157196, 
    -0.02136111, -0.02089669, -0.02097975, -0.02083927, -0.02070602, 
    -0.02048427, -0.0205206, -0.0204235, -0.02084299, -0.02056319, 
    -0.02102721, -0.02089922, -0.02193966, -0.02235028, -0.02252711, 
    -0.02268319, -0.02306753, -0.02280139, -0.02290592, -0.02265808, 
    -0.02250203, -0.02257908, -0.02210798, -0.0222899, -0.02134868, 
    -0.02174892, -0.02072152, -0.02096268, -0.02066415, -0.02081593, 
    -0.02055656, -0.02078984, -0.0203875, -0.02030096, -0.02036005, 
    -0.02013406, -0.02080285, -0.02054329, -0.02258123, -0.02256865, 
    -0.02251012, -0.02276856, -0.02278448, -0.02302424, -0.02281079, 
    -0.0227205, -0.02249303, -0.02235958, -0.02223349, -0.02195885, 
    -0.02165629, -0.0212405, -0.02094696, -0.02075255, -0.02087154, 
    -0.02076645, -0.02088396, -0.02093928, -0.02033333, -0.02067128, 
    -0.0201664, -0.02019401, -0.0204212, -0.02019089, -0.02255982, 
    -0.02263231, -0.02288585, -0.02268718, -0.02305051, -0.02284638, 
    -0.02272985, -0.02228605, -0.02218979, -0.02210088, -0.02192639, 
    -0.02170455, -0.02132101, -0.02099307, -0.0206983, -0.02071976, 
    -0.0207122, -0.02064689, -0.02080905, -0.02062039, -0.02058889, 
    -0.02067134, -0.02019771, -0.02033185, -0.02019459, -0.02028182, 
    -0.02260872, -0.02248702, -0.0225527, -0.02242935, -0.02251616, 
    -0.02213277, -0.02201915, -0.02149556, -0.02170889, -0.02137044, 
    -0.02167426, -0.02162009, -0.02135944, -0.02165774, -0.02101099, 
    -0.02144718, -0.02064435, -0.02107195, -0.02061786, -0.02069957, 
    -0.02056447, -0.02044425, -0.02029406, -0.02001992, -0.02008306, 
    -0.01985604, -0.02230686, -0.02215132, -0.02216499, -0.02200334, 
    -0.02188457, -0.02162947, -0.02122674, -0.02137727, -0.0211018, 
    -0.02104693, -0.02146579, -0.02120758, -0.02204787, -0.02190977, 
    -0.02199191, -0.02229454, -0.02134245, -0.02182564, -0.02094213, 
    -0.02119741, -0.02046134, -0.02082399, -0.0201179, -0.01982366, 
    -0.01955094, -0.01923707, -0.02206693, -0.02217208, -0.02198421, 
    -0.02172696, -0.02149115, -0.02118174, -0.02115036, -0.02109299, 
    -0.02094519, -0.02082174, -0.02107487, -0.02079091, -0.02187782, 
    -0.02130105, -0.02221194, -0.02193343, -0.02174205, -0.02182581, 
    -0.02139455, -0.02129419, -0.02089141, -0.02109864, -0.01989584, 
    -0.02041891, -0.01900169, -0.01938708, -0.02220893, -0.02206731, 
    -0.02158167, -0.02181134, -0.02116127, -0.02100436, -0.02087772, 
    -0.02071696, -0.0206997, -0.02060515, -0.02076032, -0.02061126, 
    -0.02118109, -0.02092444, -0.02163664, -0.02146099, -0.02154162, 
    -0.0216304, -0.02135759, -0.02107085, -0.02106481, -0.02097374, 
    -0.02071924, -0.02115867, -0.01982929, -0.02063956, -0.02191395, 
    -0.0216457, -0.02160772, -0.02171102, -0.02102003, -0.02126771, 
    -0.02060745, -0.02078377, -0.0204957, -0.02063832, -0.02065939, 
    -0.02084428, -0.02096026, -0.02125628, -0.02150036, -0.02169601, 
    -0.02165036, -0.02143601, -0.02105345, -0.02069812, -0.02077541, 
    -0.02051745, -0.02120771, -0.02091535, -0.02102783, -0.02073585, 
    -0.02138127, -0.02083025, -0.02152453, -0.02146271, -0.02127266, 
    -0.02089565, -0.02081324, -0.02072555, -0.02077962, -0.02104384, 
    -0.02108748, -0.02127727, -0.02132996, -0.02147616, -0.02159797, 
    -0.02148664, -0.02137036, -0.02104374, -0.02075385, -0.02044253, 
    -0.02036711, -0.02001082, -0.02030031, -0.01982486, -0.02022825, 
    -0.01953532, -0.02079883, -0.02024032, -0.02126407, -0.02115124, 
    -0.0209487, -0.02049184, -0.02073722, -0.02045057, -0.02108919, 
    -0.02142864, -0.02151744, -0.02168406, -0.02151364, -0.02152745, 
    -0.02136558, -0.02141746, -0.02103299, -0.02123861, -0.0206599, 
    -0.02045283, -0.01987969, -0.01953663, -0.01919382, -0.01904446, 
    -0.01899924, -0.01898037,
  -0.02071487, -0.02036207, -0.0204302, -0.02014902, -0.02030453, 
    -0.02012109, -0.02064288, -0.02034817, -0.02053583, -0.02068289, 
    -0.01961415, -0.02013657, -0.01908578, -0.01940857, -0.01860777, 
    -0.01913564, -0.01850308, -0.01862282, -0.0182648, -0.01836667, 
    -0.01791606, -0.01821797, -0.01768683, -0.01798773, -0.01794032, 
    -0.01822801, -0.02003038, -0.01967844, -0.02005141, -0.0200008, 
    -0.0200235, -0.0203013, -0.0204427, -0.02074211, -0.02068744, -0.0204677, 
    -0.01997808, -0.020143, -0.01972999, -0.01973922, -0.019289, -0.01949073, 
    -0.01874915, -0.01895705, -0.01836241, -0.0185102, -0.01836932, 
    -0.01841193, -0.01836877, -0.01858599, -0.01849261, -0.0186849, 
    -0.01945278, -0.01922393, -0.01991443, -0.02034128, -0.02062986, 
    -0.02083706, -0.02080764, -0.02075167, -0.02046642, -0.02020179, 
    -0.02000238, -0.01987007, -0.01974055, -0.01935347, -0.0191517, 
    -0.01870736, -0.01878683, -0.01865243, -0.01852497, -0.01831285, 
    -0.0183476, -0.01825473, -0.01865599, -0.01838834, -0.01883223, 
    -0.01870978, -0.01970536, -0.02009838, -0.02026766, -0.02041708, 
    -0.02078505, -0.02053024, -0.02063031, -0.02039304, -0.02024365, 
    -0.02031741, -0.01986646, -0.02004059, -0.01913981, -0.01952281, 
    -0.01853979, -0.01877049, -0.01848491, -0.0186301, -0.018382, 
    -0.01860514, -0.01822029, -0.01813752, -0.01819404, -0.01797791, 
    -0.01861759, -0.01836931, -0.02031947, -0.02030742, -0.0202514, 
    -0.02049881, -0.02051405, -0.0207436, -0.02053923, -0.0204528, 
    -0.02023504, -0.02010729, -0.01998659, -0.01972373, -0.01943417, 
    -0.0190363, -0.01875545, -0.01856947, -0.0186833, -0.01858277, 
    -0.01869518, -0.01874811, -0.01816848, -0.01849174, -0.01800884, 
    -0.01803524, -0.01825252, -0.01803226, -0.02029897, -0.02036837, 
    -0.0206111, -0.0204209, -0.02076876, -0.02057331, -0.02046175, 
    -0.02003691, -0.01994477, -0.01985966, -0.01969266, -0.01948035, 
    -0.01911334, -0.01879957, -0.01851758, -0.0185381, -0.01853088, 
    -0.0184684, -0.01862352, -0.01844305, -0.01841292, -0.01849179, 
    -0.01803877, -0.01816707, -0.0180358, -0.01811922, -0.02034578, 
    -0.02022928, -0.02029215, -0.02017408, -0.02025718, -0.01989019, 
    -0.01978144, -0.01928036, -0.0194845, -0.01916063, -0.01945137, 
    -0.01939953, -0.0191501, -0.01943555, -0.01881671, -0.01923406, 
    -0.01846597, -0.01887504, -0.01844063, -0.01851879, -0.01838957, 
    -0.01827457, -0.01813092, -0.01786875, -0.01792913, -0.01771205, 
    -0.02005683, -0.01990794, -0.01992103, -0.01976631, -0.01965264, 
    -0.0194085, -0.01902313, -0.01916716, -0.01890359, -0.0188511, 
    -0.01925187, -0.0190048, -0.01980893, -0.01967675, -0.01975536, 
    -0.02004503, -0.01913385, -0.01959624, -0.01875084, -0.01899507, 
    -0.01829092, -0.01863781, -0.01796245, -0.01768108, -0.01742033, 
    -0.01712028, -0.01982717, -0.01992781, -0.01974799, -0.0195018, 
    -0.01927614, -0.01898008, -0.01895005, -0.01889517, -0.01875376, 
    -0.01863566, -0.01887783, -0.01860617, -0.01964618, -0.01909423, 
    -0.01996597, -0.01969939, -0.01951624, -0.0195964, -0.0191837, 
    -0.01908768, -0.01870232, -0.01890057, -0.0177501, -0.01825034, 
    -0.0168953, -0.01726368, -0.01996309, -0.01982753, -0.01936276, 
    -0.01958255, -0.01896049, -0.01881037, -0.01868922, -0.01853543, 
    -0.01851892, -0.01842847, -0.01857691, -0.01843432, -0.01897945, 
    -0.01873391, -0.01941536, -0.01924727, -0.01932443, -0.01940939, 
    -0.01914834, -0.01887399, -0.0188682, -0.01878107, -0.01853761, 
    -0.01895801, -0.01768647, -0.01846139, -0.01968075, -0.01942404, 
    -0.01938768, -0.01948654, -0.01882537, -0.01906234, -0.01843067, 
    -0.01859934, -0.01832378, -0.0184602, -0.01848035, -0.01865723, 
    -0.01876818, -0.0190514, -0.01928495, -0.01947218, -0.01942849, 
    -0.01922338, -0.01885734, -0.01851741, -0.01859135, -0.01834458, 
    -0.01900493, -0.01872521, -0.01883283, -0.0185535, -0.019171, -0.0186438, 
    -0.01930808, -0.01924892, -0.01906707, -0.01870636, -0.01862753, 
    -0.01854365, -0.01859537, -0.01884814, -0.01888989, -0.01907148, 
    -0.0191219, -0.01926179, -0.01937835, -0.01927182, -0.01916055, 
    -0.01884805, -0.01857071, -0.01827293, -0.01820079, -0.01786005, 
    -0.0181369, -0.01768224, -0.01806799, -0.0174054, -0.01861375, 
    -0.01807953, -0.01905885, -0.01895089, -0.01875712, -0.01832009, 
    -0.0185548, -0.01828062, -0.01889153, -0.01921632, -0.01930129, 
    -0.01946074, -0.01929766, -0.01931087, -0.01915598, -0.01920563, 
    -0.01883776, -0.01903449, -0.01848085, -0.01828278, -0.01773466, 
    -0.01740665, -0.01707894, -0.01693618, -0.01689296, -0.01687492,
  -0.01736269, -0.01703655, -0.01709952, -0.01683962, -0.01698336, 
    -0.01681381, -0.01729613, -0.0170237, -0.01719717, -0.01733312, 
    -0.01634531, -0.01682811, -0.01585713, -0.01615535, -0.01541558, 
    -0.01590319, -0.0153189, -0.01542949, -0.01509884, -0.01519292, 
    -0.01477684, -0.0150556, -0.01456522, -0.01484301, -0.01479923, 
    -0.01506487, -0.01672997, -0.01640473, -0.01674941, -0.01670263, 
    -0.01672362, -0.01698037, -0.01711108, -0.01738787, -0.01733733, 
    -0.01713419, -0.01668164, -0.01683406, -0.01645236, -0.01646089, 
    -0.01604488, -0.01623127, -0.01554616, -0.01573821, -0.01518898, 
    -0.01532547, -0.01519536, -0.01523471, -0.01519485, -0.01539547, 
    -0.01530922, -0.01548682, -0.01619621, -0.01598476, -0.01662281, 
    -0.01701733, -0.0172841, -0.01747565, -0.01744845, -0.01739671, 
    -0.01713301, -0.0168884, -0.01670409, -0.01658181, -0.01646212, 
    -0.01610444, -0.01591803, -0.01550757, -0.01558097, -0.01545683, 
    -0.01533911, -0.01514321, -0.01517531, -0.01508954, -0.01546012, 
    -0.01521293, -0.01562291, -0.0155098, -0.0164296, -0.01679282, 
    -0.01694928, -0.0170874, -0.01742757, -0.017192, -0.01728451, 
    -0.01706517, -0.01692709, -0.01699526, -0.01657848, -0.0167394, 
    -0.01590704, -0.01626091, -0.0153528, -0.01556588, -0.01530212, 
    -0.01543621, -0.01520707, -0.01541316, -0.01505774, -0.01498132, 
    -0.0150335, -0.01483394, -0.01542465, -0.01519535, -0.01699717, 
    -0.01698604, -0.01693425, -0.01716295, -0.01717704, -0.01738925, 
    -0.01720032, -0.01712042, -0.01691913, -0.01680105, -0.0166895, 
    -0.01644657, -0.016179, -0.01581142, -0.01555199, -0.01538021, 
    -0.01548535, -0.01539249, -0.01549632, -0.0155452, -0.01500991, 
    -0.01530842, -0.0148625, -0.01488687, -0.01508751, -0.01488412, 
    -0.01697822, -0.01704237, -0.01726675, -0.01709093, -0.0174125, 
    -0.01723182, -0.01712869, -0.016736, -0.01665084, -0.01657219, 
    -0.01641786, -0.01622168, -0.01588259, -0.01559274, -0.01533229, 
    -0.01535124, -0.01534456, -0.01528686, -0.01543013, -0.01526345, 
    -0.01523563, -0.01530846, -0.01489014, -0.0150086, -0.01488739, 
    -0.01496442, -0.0170215, -0.01691381, -0.01697192, -0.01686278, 
    -0.0169396, -0.01660041, -0.01649991, -0.01603689, -0.01622551, 
    -0.01592628, -0.0161949, -0.016147, -0.01591655, -0.01618029, 
    -0.01560857, -0.01599412, -0.01528462, -0.01566245, -0.01526122, 
    -0.0153334, -0.01521406, -0.01510787, -0.01497522, -0.01473316, 
    -0.01478891, -0.0145885, -0.01675441, -0.01661682, -0.01662891, 
    -0.01648592, -0.01638088, -0.01615529, -0.01579925, -0.01593231, 
    -0.01568882, -0.01564034, -0.01601057, -0.01578232, -0.01652531, 
    -0.01640316, -0.01647581, -0.01674351, -0.01590153, -0.01632876, 
    -0.01554773, -0.01577333, -0.01512296, -0.01544333, -0.01481967, 
    -0.01455992, -0.01431924, -0.01404233, -0.01654217, -0.01663518, 
    -0.016469, -0.0162415, -0.016033, -0.01575948, -0.01573174, -0.01568105, 
    -0.01555042, -0.01544134, -0.01566503, -0.0154141, -0.01637491, 
    -0.01586494, -0.01667044, -0.01642408, -0.01625484, -0.01632891, 
    -0.01594759, -0.01585888, -0.01550291, -0.01568603, -0.01462363, 
    -0.01508549, -0.01383474, -0.01417466, -0.01666778, -0.0165425, 
    -0.01611302, -0.01631611, -0.01574138, -0.01560271, -0.01549081, 
    -0.01534877, -0.01533352, -0.01524999, -0.01538708, -0.01525539, 
    -0.0157589, -0.01553209, -0.01616163, -0.01600633, -0.01607761, 
    -0.01615611, -0.01591492, -0.01566148, -0.01565613, -0.01557565, 
    -0.01535078, -0.01573909, -0.01456489, -0.01528039, -0.01640685, 
    -0.01616964, -0.01613606, -0.0162274, -0.01561657, -0.01583547, 
    -0.01525202, -0.01540779, -0.01515331, -0.01527929, -0.0152979, 
    -0.01546126, -0.01556374, -0.01582537, -0.01604114, -0.01621413, 
    -0.01617376, -0.01598425, -0.0156461, -0.01533212, -0.01540041, 
    -0.01517252, -0.01578244, -0.01552406, -0.01562346, -0.01536546, 
    -0.01593585, -0.01544886, -0.0160625, -0.01600785, -0.01583984, 
    -0.01550665, -0.01543383, -0.01535636, -0.01540413, -0.0156376, 
    -0.01567617, -0.01584392, -0.0158905, -0.01601974, -0.01612743, 
    -0.016029, -0.0159262, -0.01563752, -0.01538136, -0.01510635, 
    -0.01503974, -0.01472513, -0.01498074, -0.01456098, -0.01491711, 
    -0.01430545, -0.0154211, -0.01492777, -0.01583225, -0.01573252, 
    -0.01555352, -0.01514991, -0.01536666, -0.01511345, -0.01567768, 
    -0.01597773, -0.01605623, -0.01620356, -0.01605288, -0.01606509, 
    -0.01592198, -0.01596785, -0.01562802, -0.01580975, -0.01529836, 
    -0.01511545, -0.01460938, -0.01430661, -0.01400418, -0.01387245, 
    -0.01383258, -0.01381594,
  -0.01391834, -0.01359566, -0.01365795, -0.01340094, -0.01354307, 
    -0.01337543, -0.01385247, -0.01358296, -0.01375455, -0.01388907, 
    -0.01291255, -0.01338957, -0.01243078, -0.01272501, -0.01199555, 
    -0.01247621, -0.01190033, -0.01200926, -0.01168368, -0.01177628, 
    -0.01136692, -0.01164113, -0.01115891, -0.01143199, -0.01138894, 
    -0.01165025, -0.01329255, -0.01297122, -0.01331177, -0.01326554, 
    -0.01328627, -0.01354011, -0.01366938, -0.01394326, -0.01389324, 
    -0.01369224, -0.01324479, -0.01339544, -0.01301826, -0.01302669, 
    -0.01261599, -0.01279995, -0.01212422, -0.01231351, -0.01177241, 
    -0.0119068, -0.01177869, -0.01181743, -0.01177819, -0.01197574, 
    -0.0118908, -0.01206574, -0.01276534, -0.01255667, -0.01318665, 
    -0.01357666, -0.01384056, -0.01403015, -0.01400323, -0.01395201, 
    -0.01369108, -0.01344916, -0.01326698, -0.01314615, -0.01302791, 
    -0.01267477, -0.01249085, -0.01208619, -0.01215851, -0.0120362, 
    -0.01192023, -0.01172736, -0.01175895, -0.01167453, -0.01203943, 
    -0.01179599, -0.01219985, -0.01208839, -0.01299579, -0.01335468, 
    -0.01350937, -0.01364596, -0.01398255, -0.01374944, -0.01384098, 
    -0.01362398, -0.01348742, -0.01355484, -0.01314285, -0.01330188, 
    -0.01248001, -0.01282921, -0.01193371, -0.01214364, -0.0118838, 
    -0.01201588, -0.01179022, -0.01199317, -0.01164324, -0.01156803, 
    -0.01161938, -0.01142307, -0.01200449, -0.01177868, -0.01355672, 
    -0.01354571, -0.0134945, -0.0137207, -0.01373463, -0.01394463, 
    -0.01375767, -0.01367862, -0.01347955, -0.01336281, -0.01325256, 
    -0.01301255, -0.01274836, -0.0123857, -0.01212995, -0.01196072, 
    -0.01206429, -0.01197281, -0.0120751, -0.01212327, -0.01159616, 
    -0.01189001, -0.01145115, -0.01147513, -0.01167252, -0.01147242, 
    -0.01353798, -0.01360142, -0.0138234, -0.01364945, -0.01396764, 
    -0.01378884, -0.0136868, -0.01329852, -0.01321436, -0.01313665, 
    -0.0129842, -0.01279049, -0.01245589, -0.01217011, -0.01191351, 
    -0.01193218, -0.01192561, -0.01186878, -0.01200989, -0.01184573, 
    -0.01181833, -0.01189005, -0.01147834, -0.01159488, -0.01147564, 
    -0.01155141, -0.01358078, -0.01347429, -0.01353175, -0.01342384, 
    -0.01349979, -0.01316452, -0.01306523, -0.01260811, -0.01279427, 
    -0.01249898, -0.01276405, -0.01271677, -0.01248939, -0.01274963, 
    -0.01218572, -0.01256592, -0.01186658, -0.01223883, -0.01184353, 
    -0.01191462, -0.0117971, -0.01169256, -0.01156204, -0.01132398, 
    -0.01137879, -0.01118178, -0.01331671, -0.01318073, -0.01319268, 
    -0.01305142, -0.01294767, -0.01272495, -0.01237371, -0.01250494, 
    -0.01226483, -0.01221703, -0.01258215, -0.01235701, -0.01309033, 
    -0.01296968, -0.01304143, -0.01330594, -0.01247458, -0.01289621, 
    -0.01212575, -0.01234814, -0.01170742, -0.01202289, -0.01140903, 
    -0.0111537, -0.0109173, -0.01064556, -0.01310698, -0.01319887, 
    -0.0130347, -0.01281005, -0.01260427, -0.01233449, -0.01230714, 
    -0.01225716, -0.01212841, -0.01202093, -0.01224137, -0.0119941, 
    -0.01294178, -0.01243848, -0.01323372, -0.01299034, -0.01282322, 
    -0.01289635, -0.01252001, -0.01243251, -0.01208159, -0.01226207, 
    -0.01121631, -0.01167054, -0.01044201, -0.01077538, -0.01323109, 
    -0.01310731, -0.01268324, -0.01288371, -0.01231664, -0.01217995, 
    -0.01206967, -0.01192975, -0.01191473, -0.01183247, -0.01196748, 
    -0.01183779, -0.01233392, -0.01211035, -0.01273121, -0.01257795, 
    -0.01264829, -0.01272577, -0.01248778, -0.01223787, -0.0122326, 
    -0.01215328, -0.01193173, -0.01231438, -0.01115858, -0.01186241, 
    -0.01297333, -0.01273912, -0.01270597, -0.01279613, -0.0121936, 
    -0.01240942, -0.01183448, -0.01198788, -0.01173729, -0.01186133, 
    -0.01187965, -0.01204056, -0.01214154, -0.01239946, -0.0126123, 
    -0.01278303, -0.01274318, -0.01255617, -0.01222271, -0.01191335, 
    -0.01198061, -0.0117562, -0.01235712, -0.01210243, -0.01220039, 
    -0.01194619, -0.01250843, -0.01202834, -0.01263339, -0.01257946, 
    -0.01241373, -0.01208528, -0.01201353, -0.01193722, -0.01198428, 
    -0.01221434, -0.01225235, -0.01241775, -0.01246369, -0.01259119, 
    -0.01269746, -0.01260033, -0.01249891, -0.01221425, -0.01196185, 
    -0.01169107, -0.01162552, -0.01131608, -0.01156747, -0.01115474, 
    -0.01150487, -0.01090377, -0.012001, -0.01151535, -0.01240624, 
    -0.0123079, -0.01213147, -0.01173394, -0.01194737, -0.01169806, 
    -0.01225385, -0.01254974, -0.0126272, -0.0127726, -0.01262389, 
    -0.01263594, -0.01249475, -0.01253999, -0.01220488, -0.01238405, 
    -0.01188011, -0.01170002, -0.0112023, -0.0109049, -0.01060813, 
    -0.01047897, -0.01043989, -0.01042358,
  -0.008339485, -0.008031338, -0.008090763, -0.007845741, -0.007981177, 
    -0.007821443, -0.008276523, -0.008019219, -0.008182982, -0.008311508, 
    -0.007381528, -0.007834908, -0.006925564, -0.007203795, -0.00651551, 
    -0.006968474, -0.006426045, -0.006528392, -0.006222868, -0.00630965, 
    -0.005926748, -0.006183018, -0.005732945, -0.005987479, -0.005947292, 
    -0.006191559, -0.007742555, -0.007437194, -0.007760843, -0.007716851, 
    -0.007736581, -0.007978356, -0.008101673, -0.008363315, -0.008315489, 
    -0.008123493, -0.007697113, -0.007840506, -0.007481846, -0.007489849, 
    -0.007100613, -0.007274778, -0.006636537, -0.0068149, -0.006306016, 
    -0.006432122, -0.006311907, -0.006348243, -0.006311434, -0.006496891, 
    -0.006417101, -0.006581515, -0.007241988, -0.007044517, -0.007641829, 
    -0.008013208, -0.00826514, -0.008446431, -0.008420672, -0.00837168, 
    -0.008122376, -0.007891675, -0.007718221, -0.007603323, -0.007491, 
    -0.007156229, -0.006982305, -0.006600747, -0.006668827, -0.006553722, 
    -0.006444737, -0.006263785, -0.006293396, -0.006214296, -0.006556764, 
    -0.006328127, -0.006707757, -0.006602815, -0.00746051, -0.007801689, 
    -0.007949049, -0.008079318, -0.008400895, -0.008178095, -0.008265538, 
    -0.008058346, -0.007928135, -0.007992399, -0.007600193, -0.007751431, 
    -0.006972065, -0.007302511, -0.006457401, -0.006654826, -0.006410528, 
    -0.006534619, -0.006322718, -0.00651327, -0.006184993, -0.00611462, 
    -0.006162665, -0.005979152, -0.006523913, -0.006311898, -0.007994198, 
    -0.007983697, -0.00793488, -0.008150653, -0.008163959, -0.008364623, 
    -0.008185954, -0.008110489, -0.00792063, -0.007809433, -0.007704505, 
    -0.007476424, -0.007225906, -0.006883012, -0.006641937, -0.006482769, 
    -0.006580145, -0.006494137, -0.006590317, -0.006635647, -0.006140935, 
    -0.006416354, -0.006005378, -0.006027771, -0.006212418, -0.006025246, 
    -0.007976329, -0.00803683, -0.008248743, -0.008082651, -0.008386635, 
    -0.008215724, -0.008118298, -0.007748231, -0.007668172, -0.007594294, 
    -0.007449509, -0.00726581, -0.006949277, -0.006679749, -0.006438429, 
    -0.00645596, -0.006449785, -0.006396428, -0.006528989, -0.006374796, 
    -0.006349089, -0.006416399, -0.006030772, -0.006139734, -0.006028247, 
    -0.006099071, -0.00801714, -0.007915616, -0.007970388, -0.007867552, 
    -0.007939919, -0.007620788, -0.007526448, -0.007093159, -0.007269397, 
    -0.006989989, -0.007240765, -0.007195991, -0.006980927, -0.007227104, 
    -0.00669445, -0.007053254, -0.006394358, -0.006744487, -0.006372728, 
    -0.006439463, -0.006329169, -0.006231186, -0.006109014, -0.005886694, 
    -0.005937819, -0.005754232, -0.00776555, -0.0076362, -0.007647562, 
    -0.007513327, -0.007414846, -0.007203738, -0.006871688, -0.006995616, 
    -0.006768991, -0.006723947, -0.007068601, -0.006855929, -0.007550284, 
    -0.00743573, -0.00750384, -0.007755293, -0.006966931, -0.007366025, 
    -0.006637986, -0.006847566, -0.006245107, -0.006541212, -0.005966051, 
    -0.005728099, -0.005508538, -0.005257097, -0.007566108, -0.007653449, 
    -0.007497451, -0.007284348, -0.007089523, -0.006834684, -0.00680889, 
    -0.006761763, -0.006640487, -0.006539369, -0.006746878, -0.006514145, 
    -0.007409254, -0.006932838, -0.007686589, -0.007455339, -0.00729683, 
    -0.007366165, -0.007009857, -0.006927196, -0.006596422, -0.006766398, 
    -0.005786373, -0.006210561, -0.00506946, -0.005377094, -0.007684085, 
    -0.007566418, -0.007164247, -0.007354179, -0.006817852, -0.006689012, 
    -0.006585208, -0.006453676, -0.006439569, -0.006362353, -0.006489128, 
    -0.006367344, -0.006834147, -0.006623485, -0.007209663, -0.007064637, 
    -0.007131172, -0.00720451, -0.006979408, -0.006743581, -0.006738618, 
    -0.006663895, -0.00645554, -0.006815722, -0.005732642, -0.00639045, 
    -0.00743919, -0.007217156, -0.007185765, -0.007271161, -0.006701871, 
    -0.006905398, -0.006364233, -0.006508301, -0.0062731, -0.006389432, 
    -0.006406636, -0.006557827, -0.006652844, -0.006895993, -0.007097124, 
    -0.007258747, -0.007221001, -0.007044042, -0.006729297, -0.006438279, 
    -0.006501469, -0.006290823, -0.006856039, -0.006616032, -0.006708271, 
    -0.006469118, -0.006998918, -0.006546338, -0.007117067, -0.00706606, 
    -0.00690947, -0.00659989, -0.006532414, -0.006460697, -0.00650491, 
    -0.006721408, -0.006757232, -0.006913262, -0.006956647, -0.007077151, 
    -0.007177708, -0.007085797, -0.006989923, -0.006721328, -0.006483831, 
    -0.006229792, -0.006168406, -0.005879333, -0.006114092, -0.005729071, 
    -0.006055566, -0.005495992, -0.006520627, -0.006065362, -0.006902398, 
    -0.006809608, -0.006643365, -0.006269957, -0.006470233, -0.006236337, 
    -0.00675864, -0.007037962, -0.007111213, -0.007248861, -0.007108083, 
    -0.007119481, -0.006985988, -0.007028746, -0.006712503, -0.006881453, 
    -0.006407061, -0.006238176, -0.00577333, -0.005497045, -0.005222553, 
    -0.005103489, -0.00506751, -0.005052504,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  439.2171, 440.8315, 440.5177, 441.8204, 441.0974, 441.9509, 439.5443, 
    440.8958, 440.0334, 439.3623, 444.3556, 441.8785, 446.9357, 445.3498, 
    449.3393, 446.6889, 449.8748, 449.2623, 451.1061, 450.5774, 452.9413, 
    451.3502, 454.1688, 452.5608, 452.8123, 451.2979, 442.376, 444.0469, 
    442.2772, 442.5152, 442.4083, 441.1124, 440.4604, 439.0935, 439.3416, 
    440.3455, 442.6223, 441.8484, 443.7995, 443.7554, 445.9337, 444.9508, 
    448.6211, 447.576, 450.5995, 449.8381, 450.5638, 450.3436, 450.5667, 
    449.4502, 449.9284, 448.9466, 445.1349, 446.2532, 442.9227, 440.9278, 
    439.6037, 438.6644, 438.7971, 439.0503, 440.3514, 441.5742, 442.5077, 
    443.1327, 443.7491, 445.6188, 446.6094, 448.8328, 448.4307, 449.1117, 
    449.7624, 450.8564, 450.6762, 451.1586, 449.0935, 450.4655, 448.2019, 
    448.8204, 443.918, 442.057, 441.2685, 440.578, 438.8992, 440.0591, 
    439.6017, 440.6886, 441.3796, 441.0377, 443.1498, 442.328, 446.6682, 
    444.7956, 449.6864, 448.5132, 449.9679, 449.2252, 450.4983, 449.3524, 
    451.3382, 451.7714, 451.4753, 452.6127, 449.289, 450.5639, 441.0282, 
    441.084, 441.3436, 440.2029, 440.1331, 439.0868, 440.0178, 440.4138, 
    441.4196, 442.0154, 442.582, 443.8295, 445.2254, 447.1812, 448.5892, 
    449.5345, 448.9547, 449.4666, 448.8944, 448.6263, 451.6091, 449.9329, 
    452.449, 452.3095, 451.1702, 452.3252, 441.1231, 440.8023, 439.6892, 
    440.5604, 438.9729, 439.8619, 440.3729, 442.3455, 442.7793, 443.1821, 
    443.9781, 445.0011, 446.799, 448.3666, 449.8002, 449.695, 449.7321, 
    450.0528, 449.2587, 450.1832, 450.3386, 449.9326, 452.2908, 451.6164, 
    452.3065, 451.8673, 440.9065, 441.4464, 441.1546, 441.7034, 441.3168, 
    443.0376, 443.5542, 445.9763, 444.981, 446.5652, 445.1417, 445.3938, 
    446.6175, 445.2184, 448.2803, 446.2036, 450.0652, 447.9872, 450.1957, 
    449.794, 450.459, 451.0553, 451.8059, 453.193, 452.8715, 454.0327, 
    442.2518, 442.9534, 442.8914, 443.6262, 444.1701, 445.35, 447.2466, 
    446.5328, 447.8435, 448.107, 446.1158, 447.338, 443.4232, 444.0546, 
    443.6784, 442.3072, 446.6976, 444.4414, 448.6126, 447.3864, 450.9703, 
    449.1862, 452.6947, 454.1999, 455.618, 457.2798, 443.3364, 442.8593, 
    443.7135, 444.8974, 445.9967, 447.4612, 447.611, 447.8858, 448.5977, 
    449.1969, 447.973, 449.3472, 444.2016, 446.8936, 442.6793, 443.9462, 
    444.8274, 444.4405, 446.4512, 446.926, 448.8584, 447.8587, 453.8284, 
    451.1817, 458.5464, 456.4817, 442.6928, 443.3346, 445.5731, 444.5072, 
    447.5589, 448.312, 448.9247, 449.7088, 449.7934, 450.2584, 449.4965, 
    450.2281, 447.4643, 448.6982, 445.3166, 446.1384, 445.7602, 445.3456, 
    446.6257, 447.9923, 448.0211, 448.4599, 449.6984, 447.5713, 454.1714, 
    450.0894, 444.0352, 445.2747, 445.4514, 444.971, 448.2365, 447.0518, 
    450.247, 449.382, 450.7996, 450.0949, 449.9913, 449.0872, 448.5249, 
    447.1061, 445.9536, 445.0406, 445.2528, 446.2559, 448.0758, 449.8012, 
    449.423, 450.6918, 447.3372, 448.7423, 448.1991, 449.6162, 446.5139, 
    449.1562, 445.8402, 446.1302, 447.0283, 448.838, 449.2383, 449.6667, 
    449.4023, 448.122, 447.9123, 447.0063, 446.7566, 446.067, 445.4969, 
    446.0179, 446.5656, 448.1224, 449.5283, 451.0639, 451.44, 453.2398, 
    451.7749, 454.1942, 452.1377, 455.7006, 449.309, 452.0765, 447.069, 
    447.6068, 448.581, 450.819, 449.6096, 451.024, 447.9041, 446.2907, 
    445.8734, 445.0962, 445.8912, 445.8265, 446.588, 446.3431, 448.1741, 
    447.1901, 449.9888, 451.0128, 453.9111, 455.6933, 457.5109, 458.3148, 
    458.5596, 458.662 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  7.623549e-08, 7.644416e-08, 7.640361e-08, 7.657187e-08, 7.647855e-08, 
    7.658871e-08, 7.627782e-08, 7.645243e-08, 7.634097e-08, 7.62543e-08, 
    7.689825e-08, 7.657938e-08, 7.722948e-08, 7.702619e-08, 7.75368e-08, 
    7.719783e-08, 7.760514e-08, 7.752706e-08, 7.776212e-08, 7.769479e-08, 
    7.79953e-08, 7.77932e-08, 7.815109e-08, 7.794706e-08, 7.797897e-08, 
    7.778652e-08, 7.664359e-08, 7.685854e-08, 7.663084e-08, 7.66615e-08, 
    7.664775e-08, 7.648046e-08, 7.639613e-08, 7.621956e-08, 7.625163e-08, 
    7.638132e-08, 7.667528e-08, 7.657553e-08, 7.682698e-08, 7.682131e-08, 
    7.710113e-08, 7.697498e-08, 7.744517e-08, 7.731157e-08, 7.76976e-08, 
    7.760053e-08, 7.769304e-08, 7.766499e-08, 7.76934e-08, 7.755104e-08, 
    7.761204e-08, 7.748676e-08, 7.69986e-08, 7.714208e-08, 7.671404e-08, 
    7.64565e-08, 7.628547e-08, 7.616406e-08, 7.618123e-08, 7.621394e-08, 
    7.638208e-08, 7.654015e-08, 7.666058e-08, 7.674113e-08, 7.682049e-08, 
    7.706056e-08, 7.718769e-08, 7.747217e-08, 7.742086e-08, 7.750779e-08, 
    7.759088e-08, 7.773031e-08, 7.770736e-08, 7.776877e-08, 7.750553e-08, 
    7.768048e-08, 7.739163e-08, 7.747064e-08, 7.684195e-08, 7.660245e-08, 
    7.650053e-08, 7.64114e-08, 7.619442e-08, 7.634426e-08, 7.62852e-08, 
    7.642574e-08, 7.651501e-08, 7.647086e-08, 7.674333e-08, 7.663741e-08, 
    7.719521e-08, 7.6955e-08, 7.758118e-08, 7.743139e-08, 7.761709e-08, 
    7.752234e-08, 7.768467e-08, 7.753858e-08, 7.779164e-08, 7.784672e-08, 
    7.780908e-08, 7.79537e-08, 7.753048e-08, 7.769302e-08, 7.646963e-08, 
    7.647682e-08, 7.651037e-08, 7.636287e-08, 7.635385e-08, 7.621868e-08, 
    7.633896e-08, 7.639017e-08, 7.652019e-08, 7.659708e-08, 7.667015e-08, 
    7.683081e-08, 7.701018e-08, 7.726096e-08, 7.744111e-08, 7.756182e-08, 
    7.748781e-08, 7.755315e-08, 7.74801e-08, 7.744587e-08, 7.782607e-08, 
    7.76126e-08, 7.79329e-08, 7.791519e-08, 7.777024e-08, 7.791719e-08, 
    7.648188e-08, 7.644044e-08, 7.629653e-08, 7.640916e-08, 7.620396e-08, 
    7.631881e-08, 7.638484e-08, 7.66396e-08, 7.669559e-08, 7.674747e-08, 
    7.684995e-08, 7.698143e-08, 7.721203e-08, 7.741262e-08, 7.759571e-08, 
    7.75823e-08, 7.758702e-08, 7.762791e-08, 7.752661e-08, 7.764454e-08, 
    7.766432e-08, 7.761258e-08, 7.791282e-08, 7.782705e-08, 7.791481e-08, 
    7.785898e-08, 7.645392e-08, 7.652364e-08, 7.648596e-08, 7.65568e-08, 
    7.650689e-08, 7.672879e-08, 7.679531e-08, 7.710651e-08, 7.697884e-08, 
    7.718206e-08, 7.699949e-08, 7.703184e-08, 7.718864e-08, 7.700937e-08, 
    7.740154e-08, 7.713565e-08, 7.762949e-08, 7.7364e-08, 7.764613e-08, 
    7.759493e-08, 7.767972e-08, 7.775563e-08, 7.785115e-08, 7.802734e-08, 
    7.798656e-08, 7.813389e-08, 7.662758e-08, 7.671798e-08, 7.671004e-08, 
    7.680465e-08, 7.687462e-08, 7.702625e-08, 7.726938e-08, 7.717797e-08, 
    7.73458e-08, 7.737948e-08, 7.712452e-08, 7.728104e-08, 7.67785e-08, 
    7.685969e-08, 7.681136e-08, 7.663471e-08, 7.7199e-08, 7.690944e-08, 
    7.744408e-08, 7.728728e-08, 7.774481e-08, 7.751729e-08, 7.79641e-08, 
    7.815497e-08, 7.833466e-08, 7.85445e-08, 7.676734e-08, 7.670592e-08, 
    7.681592e-08, 7.696804e-08, 7.710922e-08, 7.729684e-08, 7.731605e-08, 
    7.735118e-08, 7.744221e-08, 7.751873e-08, 7.736227e-08, 7.753791e-08, 
    7.687849e-08, 7.722414e-08, 7.668267e-08, 7.684573e-08, 7.695908e-08, 
    7.690938e-08, 7.716753e-08, 7.722835e-08, 7.747545e-08, 7.734774e-08, 
    7.810785e-08, 7.777165e-08, 7.87043e-08, 7.844376e-08, 7.668445e-08, 
    7.676714e-08, 7.705483e-08, 7.691796e-08, 7.730937e-08, 7.740568e-08, 
    7.748397e-08, 7.758402e-08, 7.759483e-08, 7.765411e-08, 7.755698e-08, 
    7.765028e-08, 7.729724e-08, 7.745503e-08, 7.702198e-08, 7.712739e-08, 
    7.70789e-08, 7.70257e-08, 7.718989e-08, 7.736472e-08, 7.73685e-08, 
    7.742454e-08, 7.758241e-08, 7.731096e-08, 7.815116e-08, 7.763233e-08, 
    7.68573e-08, 7.701648e-08, 7.703925e-08, 7.697759e-08, 7.739602e-08, 
    7.724444e-08, 7.765266e-08, 7.754237e-08, 7.772309e-08, 7.763329e-08, 
    7.762007e-08, 7.750472e-08, 7.743289e-08, 7.725138e-08, 7.710367e-08, 
    7.698654e-08, 7.701378e-08, 7.714245e-08, 7.737543e-08, 7.75958e-08, 
    7.754753e-08, 7.770936e-08, 7.7281e-08, 7.746063e-08, 7.73912e-08, 
    7.757223e-08, 7.717554e-08, 7.751326e-08, 7.708917e-08, 7.712637e-08, 
    7.724142e-08, 7.747279e-08, 7.752402e-08, 7.757865e-08, 7.754495e-08, 
    7.738135e-08, 7.735456e-08, 7.723864e-08, 7.720661e-08, 7.711827e-08, 
    7.704512e-08, 7.711195e-08, 7.718212e-08, 7.738143e-08, 7.756099e-08, 
    7.77567e-08, 7.780461e-08, 7.803313e-08, 7.784707e-08, 7.815405e-08, 
    7.7893e-08, 7.834487e-08, 7.753288e-08, 7.788538e-08, 7.724667e-08, 
    7.731551e-08, 7.743999e-08, 7.772545e-08, 7.757139e-08, 7.775158e-08, 
    7.735351e-08, 7.714686e-08, 7.709342e-08, 7.699366e-08, 7.709571e-08, 
    7.708741e-08, 7.718505e-08, 7.715368e-08, 7.738805e-08, 7.726216e-08, 
    7.761973e-08, 7.775017e-08, 7.811844e-08, 7.834409e-08, 7.857378e-08, 
    7.867516e-08, 7.8706e-08, 7.871891e-08 ;

 SOM_C_LEACHED =
  2.809888e-20, 1.821581e-20, 6.040847e-21, -7.491634e-22, -7.922864e-21, 
    3.951862e-21, -4.114505e-20, 1.418723e-20, -2.27792e-20, -7.763929e-21, 
    1.765267e-20, -4.259754e-20, -3.398543e-20, 9.341675e-22, 2.027686e-20, 
    -2.493581e-21, -1.47718e-20, 7.729735e-20, -7.42878e-21, -3.809609e-20, 
    1.184947e-20, 2.867801e-20, 1.463607e-20, -2.169957e-20, 2.162908e-21, 
    -5.433796e-20, 5.979293e-20, -3.414519e-20, -1.024302e-20, -1.962833e-20, 
    9.963626e-21, -2.163411e-20, -1.280956e-21, 1.118988e-20, -1.295861e-20, 
    4.70269e-20, -3.184382e-20, 8.797483e-20, 3.451883e-20, 2.228501e-20, 
    -6.941891e-21, 3.920831e-20, -6.494948e-20, 4.62841e-20, 1.817002e-20, 
    2.025187e-20, 2.039864e-20, 5.486891e-20, 2.619333e-20, 5.744685e-20, 
    7.391042e-21, -4.101829e-20, -7.241622e-21, 3.548757e-20, -1.599002e-20, 
    1.317372e-20, 2.476363e-20, 4.997515e-20, -1.071016e-20, 4.722794e-20, 
    5.189383e-21, 3.890948e-20, -5.294484e-20, 5.787946e-20, -1.22386e-20, 
    -6.004579e-21, 1.03429e-20, 3.105455e-20, -2.833828e-20, -1.176159e-20, 
    2.040698e-20, -2.059033e-20, 6.393345e-20, -8.22147e-20, 2.297399e-20, 
    -8.283076e-21, -2.208824e-20, -3.63893e-20, -1.122368e-20, -1.852241e-20, 
    -1.197239e-20, -1.845174e-20, -6.608003e-20, -4.408897e-20, 2.919826e-20, 
    -4.990708e-20, -4.239545e-20, -1.964464e-20, 1.186066e-20, -3.442427e-20, 
    3.457026e-20, -4.609147e-20, -4.10366e-20, 4.408782e-21, 2.592682e-21, 
    5.046521e-20, 8.277598e-21, -6.569646e-21, -5.341622e-20, -6.088624e-21, 
    -5.450454e-20, -1.510534e-20, 3.232505e-20, 1.891492e-20, 3.296493e-20, 
    2.067808e-20, -5.944884e-21, 4.0583e-21, -1.410046e-20, 5.901578e-20, 
    1.014921e-20, 7.150936e-20, -4.002061e-20, -1.894064e-20, -1.76268e-20, 
    -4.609947e-21, -3.406753e-20, -6.012908e-20, -1.476276e-20, 4.067673e-20, 
    4.151403e-20, 2.323532e-20, -2.741435e-21, -2.344514e-20, -4.47556e-20, 
    -4.363948e-20, -3.415481e-20, 2.253173e-20, 1.787976e-20, 4.13025e-22, 
    -5.282238e-21, 3.981681e-20, -8.912677e-20, -4.0854e-20, 8.461527e-21, 
    -2.01787e-21, 8.738355e-21, 5.39051e-20, -3.500949e-20, 5.676003e-20, 
    -8.705597e-21, -4.608622e-20, 2.033882e-20, -8.705164e-20, -9.09775e-21, 
    1.311701e-20, 7.554779e-21, 4.740618e-20, -4.664798e-20, 8.45854e-21, 
    7.340741e-20, -4.841961e-20, 1.779544e-20, -3.508578e-20, -4.386603e-20, 
    -6.658364e-21, 7.155478e-20, -1.279828e-20, -2.913863e-20, -1.188797e-20, 
    -3.514935e-20, -1.267373e-20, -8.670112e-20, -4.517238e-20, 2.483796e-20, 
    -7.806586e-20, 3.217869e-20, -5.714686e-20, -9.262547e-20, -2.466372e-20, 
    1.545674e-21, -6.388395e-20, -3.549986e-20, -1.01364e-21, 8.598193e-20, 
    2.348098e-20, 1.710361e-20, 9.075204e-21, 3.273242e-20, -3.81011e-20, 
    -4.742997e-21, 3.3278e-20, -1.932172e-20, -2.972324e-20, -6.974706e-20, 
    -2.055161e-20, -3.057654e-20, 1.7111e-20, 2.38431e-20, 2.146261e-20, 
    2.393656e-20, 5.128911e-20, 4.078845e-21, -1.503574e-20, -2.014619e-20, 
    6.324673e-20, -3.29244e-20, -6.596495e-20, -3.543289e-20, 9.771485e-21, 
    -1.624688e-20, -1.051814e-20, 2.99719e-20, -1.592346e-21, 2.373231e-20, 
    -5.079711e-20, 3.114706e-20, 1.802022e-20, -4.023559e-20, 9.059299e-20, 
    -1.529744e-20, 1.309021e-20, 1.12145e-19, 1.08217e-20, 3.780259e-20, 
    -1.022362e-19, -3.597768e-20, 3.406517e-20, 4.829199e-20, 7.012913e-21, 
    7.809338e-20, -1.22136e-20, -4.092412e-20, 4.517818e-20, -2.37817e-20, 
    2.324903e-20, -6.100437e-20, 4.920758e-21, 3.118122e-20, 3.930027e-20, 
    -2.329646e-20, 5.449758e-20, -3.006602e-20, 4.089939e-20, -4.24941e-20, 
    1.120702e-20, -1.153395e-20, -5.285337e-20, -6.43443e-21, 2.000526e-20, 
    3.150967e-20, -2.470856e-20, -1.73497e-20, -2.356424e-20, -5.386705e-20, 
    1.720688e-20, 7.370461e-20, -1.70804e-23, -3.895697e-20, 7.977052e-20, 
    7.834064e-21, 4.937019e-21, -2.433862e-20, -4.158331e-20, 1.117846e-20, 
    2.015362e-20, 4.416384e-20, 1.088941e-20, 3.956723e-20, -1.46257e-20, 
    9.128197e-21, 2.280497e-20, 3.096252e-20, 2.438317e-20, -2.33172e-20, 
    3.021856e-20, -7.697426e-20, -4.91419e-21, -5.475145e-20, 2.239612e-20, 
    2.383523e-20, 5.656524e-20, 1.23527e-20, -1.492084e-20, 1.256636e-20, 
    -3.62617e-20, -6.317236e-20, 1.982102e-20, 6.057241e-20, 3.354602e-20, 
    4.489986e-20, -4.663711e-20, -1.891407e-20, -3.322351e-20, -6.346472e-20, 
    1.872986e-20, 3.797425e-20, 3.826811e-20, -6.134148e-21, -3.502809e-20, 
    -1.122913e-21, 3.361864e-21, 1.068336e-20, 1.472259e-20, 7.586608e-20, 
    1.287718e-20, -3.624462e-21, -2.179232e-20, 4.081502e-20, -1.83366e-20, 
    -4.285495e-20, 1.074181e-20, 3.209785e-20, -5.221828e-21, 6.062772e-21, 
    5.867871e-20, 2.00472e-20, 8.075593e-22, -9.30256e-20, -8.806883e-21, 
    3.506715e-20, -2.021627e-20, 6.053281e-21, -9.169035e-20, 4.241523e-20, 
    5.845692e-20, 5.890741e-21, -9.230848e-21, -1.724104e-20, 3.593698e-20, 
    -5.771154e-20, -2.64342e-20, 2.757362e-20, -3.418338e-20, 2.615469e-20, 
    -1.062223e-20, -2.867244e-20, -5.697314e-21, -5.45288e-20, 3.385665e-20, 
    -8.477991e-21, -2.916945e-20, 9.900143e-20, 5.20836e-20, 9.107257e-21, 
    2.301682e-20, -1.090054e-20, 5.03339e-20 ;

 SR =
  7.623649e-08, 7.644516e-08, 7.640461e-08, 7.657286e-08, 7.647954e-08, 
    7.658971e-08, 7.627882e-08, 7.645342e-08, 7.634197e-08, 7.62553e-08, 
    7.689925e-08, 7.658038e-08, 7.723048e-08, 7.70272e-08, 7.753781e-08, 
    7.719884e-08, 7.760615e-08, 7.752807e-08, 7.776314e-08, 7.76958e-08, 
    7.799632e-08, 7.779421e-08, 7.815211e-08, 7.794808e-08, 7.797998e-08, 
    7.778754e-08, 7.664459e-08, 7.685954e-08, 7.663184e-08, 7.66625e-08, 
    7.664875e-08, 7.648146e-08, 7.639712e-08, 7.622056e-08, 7.625263e-08, 
    7.638231e-08, 7.667629e-08, 7.657653e-08, 7.682798e-08, 7.682231e-08, 
    7.710213e-08, 7.697598e-08, 7.744618e-08, 7.731258e-08, 7.769862e-08, 
    7.760154e-08, 7.769405e-08, 7.766601e-08, 7.769442e-08, 7.755205e-08, 
    7.761304e-08, 7.748777e-08, 7.69996e-08, 7.714308e-08, 7.671504e-08, 
    7.64575e-08, 7.628647e-08, 7.616506e-08, 7.618222e-08, 7.621494e-08, 
    7.638307e-08, 7.654115e-08, 7.666159e-08, 7.674213e-08, 7.682149e-08, 
    7.706157e-08, 7.718869e-08, 7.747317e-08, 7.742187e-08, 7.750881e-08, 
    7.759189e-08, 7.773131e-08, 7.770838e-08, 7.776979e-08, 7.750653e-08, 
    7.768149e-08, 7.739264e-08, 7.747165e-08, 7.684295e-08, 7.660345e-08, 
    7.650154e-08, 7.64124e-08, 7.619542e-08, 7.634526e-08, 7.628619e-08, 
    7.642673e-08, 7.651601e-08, 7.647186e-08, 7.674434e-08, 7.663841e-08, 
    7.719622e-08, 7.695601e-08, 7.758219e-08, 7.74324e-08, 7.76181e-08, 
    7.752336e-08, 7.768568e-08, 7.75396e-08, 7.779266e-08, 7.784774e-08, 
    7.781009e-08, 7.795472e-08, 7.753149e-08, 7.769404e-08, 7.647062e-08, 
    7.647782e-08, 7.651137e-08, 7.636387e-08, 7.635484e-08, 7.621968e-08, 
    7.633997e-08, 7.639117e-08, 7.65212e-08, 7.659807e-08, 7.667116e-08, 
    7.683181e-08, 7.701119e-08, 7.726197e-08, 7.744212e-08, 7.756284e-08, 
    7.748882e-08, 7.755416e-08, 7.748111e-08, 7.744688e-08, 7.782709e-08, 
    7.761361e-08, 7.793392e-08, 7.791621e-08, 7.777125e-08, 7.791819e-08, 
    7.648288e-08, 7.644144e-08, 7.629752e-08, 7.641015e-08, 7.620496e-08, 
    7.631981e-08, 7.638584e-08, 7.66406e-08, 7.669659e-08, 7.674847e-08, 
    7.685095e-08, 7.698243e-08, 7.721304e-08, 7.741363e-08, 7.759672e-08, 
    7.758331e-08, 7.758803e-08, 7.762892e-08, 7.752763e-08, 7.764555e-08, 
    7.766533e-08, 7.76136e-08, 7.791383e-08, 7.782807e-08, 7.791583e-08, 
    7.785999e-08, 7.645492e-08, 7.652464e-08, 7.648696e-08, 7.65578e-08, 
    7.650789e-08, 7.672979e-08, 7.679631e-08, 7.710752e-08, 7.697984e-08, 
    7.718307e-08, 7.700049e-08, 7.703284e-08, 7.718965e-08, 7.701037e-08, 
    7.740255e-08, 7.713665e-08, 7.76305e-08, 7.736501e-08, 7.764714e-08, 
    7.759594e-08, 7.768072e-08, 7.775665e-08, 7.785217e-08, 7.802836e-08, 
    7.798757e-08, 7.813491e-08, 7.662858e-08, 7.671898e-08, 7.671105e-08, 
    7.680566e-08, 7.687562e-08, 7.702726e-08, 7.727039e-08, 7.717897e-08, 
    7.73468e-08, 7.738048e-08, 7.712552e-08, 7.728205e-08, 7.67795e-08, 
    7.686069e-08, 7.681236e-08, 7.66357e-08, 7.720001e-08, 7.691045e-08, 
    7.744509e-08, 7.728828e-08, 7.774582e-08, 7.751829e-08, 7.796511e-08, 
    7.815598e-08, 7.833569e-08, 7.854553e-08, 7.676834e-08, 7.670692e-08, 
    7.681692e-08, 7.696904e-08, 7.711023e-08, 7.729785e-08, 7.731705e-08, 
    7.735219e-08, 7.744323e-08, 7.751974e-08, 7.736328e-08, 7.753892e-08, 
    7.687949e-08, 7.722515e-08, 7.668368e-08, 7.684673e-08, 7.696008e-08, 
    7.691038e-08, 7.716854e-08, 7.722935e-08, 7.747646e-08, 7.734874e-08, 
    7.810886e-08, 7.777265e-08, 7.870533e-08, 7.844478e-08, 7.668545e-08, 
    7.676814e-08, 7.705584e-08, 7.691897e-08, 7.731038e-08, 7.740669e-08, 
    7.748498e-08, 7.758503e-08, 7.759585e-08, 7.765512e-08, 7.755798e-08, 
    7.765129e-08, 7.729825e-08, 7.745604e-08, 7.702298e-08, 7.71284e-08, 
    7.707991e-08, 7.702671e-08, 7.71909e-08, 7.736573e-08, 7.736951e-08, 
    7.742555e-08, 7.758342e-08, 7.731197e-08, 7.815218e-08, 7.763335e-08, 
    7.68583e-08, 7.701748e-08, 7.704026e-08, 7.697859e-08, 7.739703e-08, 
    7.724544e-08, 7.765367e-08, 7.754338e-08, 7.77241e-08, 7.76343e-08, 
    7.762108e-08, 7.750573e-08, 7.74339e-08, 7.725239e-08, 7.710467e-08, 
    7.698755e-08, 7.701478e-08, 7.714345e-08, 7.737644e-08, 7.759681e-08, 
    7.754854e-08, 7.771037e-08, 7.728201e-08, 7.746164e-08, 7.739221e-08, 
    7.757325e-08, 7.717654e-08, 7.751427e-08, 7.709018e-08, 7.712737e-08, 
    7.724243e-08, 7.74738e-08, 7.752503e-08, 7.757966e-08, 7.754596e-08, 
    7.738236e-08, 7.735557e-08, 7.723964e-08, 7.720762e-08, 7.711928e-08, 
    7.704612e-08, 7.711296e-08, 7.718313e-08, 7.738244e-08, 7.7562e-08, 
    7.775772e-08, 7.780563e-08, 7.803415e-08, 7.784809e-08, 7.815506e-08, 
    7.789401e-08, 7.834588e-08, 7.753389e-08, 7.788639e-08, 7.724768e-08, 
    7.731652e-08, 7.744099e-08, 7.772646e-08, 7.757239e-08, 7.775259e-08, 
    7.735452e-08, 7.714787e-08, 7.709443e-08, 7.699466e-08, 7.709671e-08, 
    7.708842e-08, 7.718606e-08, 7.715469e-08, 7.738906e-08, 7.726317e-08, 
    7.762075e-08, 7.775118e-08, 7.811946e-08, 7.834512e-08, 7.857481e-08, 
    7.867618e-08, 7.870703e-08, 7.871993e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.341361, -0.3413828, -0.3413818, -0.3413859, -0.3413837, -0.3413863, 
    -0.3413621, -0.3413829, -0.3413637, -0.3413616, -0.3413936, -0.3413861, 
    -0.3414276, -0.341397, -0.3414353, -0.3414268, -0.3414371, -0.3414352, 
    -0.3414412, -0.3414395, -0.3414468, -0.3414419, -0.3414508, -0.3414457, 
    -0.3414465, -0.3414418, -0.3413877, -0.3413927, -0.3413874, -0.3413881, 
    -0.3413878, -0.3413837, -0.3413815, -0.3413607, -0.3413615, -0.3413812, 
    -0.3413884, -0.341386, -0.3413922, -0.3413921, -0.3413989, -0.3413958, 
    -0.3414331, -0.3414298, -0.3414395, -0.3414371, -0.3414394, -0.3414387, 
    -0.3414394, -0.3414358, -0.3414373, -0.3414342, -0.3413964, -0.3414255, 
    -0.3413894, -0.3413829, -0.3413623, -0.3413594, -0.3413598, -0.3413605, 
    -0.3413812, -0.3413852, -0.3413882, -0.3413901, -0.3413921, -0.3413977, 
    -0.3414266, -0.3414338, -0.3414326, -0.3414347, -0.3414368, -0.3414403, 
    -0.3414398, -0.3414413, -0.3414347, -0.341439, -0.3414319, -0.3414338, 
    -0.3413922, -0.3413867, -0.341384, -0.341382, -0.3413601, -0.3413637, 
    -0.3413623, -0.3413824, -0.3413846, -0.3413835, -0.3413902, -0.3413876, 
    -0.3414268, -0.3413953, -0.3414366, -0.3414328, -0.3414375, -0.3414351, 
    -0.3414392, -0.3414355, -0.3414419, -0.3414432, -0.3414423, -0.341446, 
    -0.3414353, -0.3414394, -0.3413835, -0.3413836, -0.3413845, -0.3413807, 
    -0.341364, -0.3413607, -0.3413636, -0.3413815, -0.3413847, -0.3413866, 
    -0.3413883, -0.3413923, -0.3413966, -0.3414285, -0.341433, -0.3414361, 
    -0.3414343, -0.3414359, -0.3414341, -0.3414332, -0.3414427, -0.3414373, 
    -0.3414454, -0.341445, -0.3414413, -0.341445, -0.3413838, -0.3413827, 
    -0.3413626, -0.341382, -0.3413603, -0.3413631, -0.3413813, -0.3413875, 
    -0.341389, -0.3413903, -0.3413928, -0.341396, -0.3414272, -0.3414323, 
    -0.341437, -0.3414367, -0.3414367, -0.3414378, -0.3414352, -0.3414382, 
    -0.3414387, -0.3414374, -0.3414449, -0.3414428, -0.341445, -0.3414436, 
    -0.3413831, -0.3413848, -0.3413838, -0.3413856, -0.3413843, -0.3413897, 
    -0.3413913, -0.3413989, -0.3413959, -0.3414265, -0.3413964, -0.3413972, 
    -0.3414265, -0.3413967, -0.3414319, -0.3414252, -0.3414378, -0.3414309, 
    -0.3414382, -0.341437, -0.3414391, -0.3414409, -0.3414434, -0.3414477, 
    -0.3414467, -0.3414504, -0.3413873, -0.3413895, -0.3413894, -0.3413917, 
    -0.3413934, -0.3413971, -0.3414287, -0.3414265, -0.3414307, -0.3414315, 
    -0.3414251, -0.341429, -0.341391, -0.3413929, -0.3413918, -0.3413875, 
    -0.3414269, -0.3413941, -0.3414331, -0.3414292, -0.3414407, -0.3414349, 
    -0.3414462, -0.3414508, -0.3414555, -0.3414606, -0.3413907, -0.3413893, 
    -0.341392, -0.3413956, -0.3414247, -0.3414294, -0.3414299, -0.3414308, 
    -0.3414331, -0.341435, -0.341431, -0.3414355, -0.3413932, -0.3414275, 
    -0.3413886, -0.3413925, -0.3413954, -0.3413942, -0.3414262, -0.3414277, 
    -0.3414339, -0.3414307, -0.3414496, -0.3414412, -0.3414647, -0.3414581, 
    -0.3413887, -0.3413908, -0.3413977, -0.3413944, -0.3414298, -0.3414322, 
    -0.3414342, -0.3414366, -0.341437, -0.3414384, -0.341436, -0.3414383, 
    -0.3414294, -0.3414334, -0.341397, -0.3414252, -0.3413984, -0.3413971, 
    -0.3414268, -0.3414311, -0.3414313, -0.3414326, -0.3414362, -0.3414298, 
    -0.3414505, -0.3414375, -0.341393, -0.3413967, -0.3413974, -0.3413959, 
    -0.3414319, -0.3414281, -0.3414384, -0.3414356, -0.3414402, -0.3414379, 
    -0.3414376, -0.3414347, -0.3414329, -0.3414283, -0.341399, -0.3413962, 
    -0.3413968, -0.3414255, -0.3414313, -0.3414369, -0.3414357, -0.3414398, 
    -0.3414291, -0.3414335, -0.3414317, -0.3414364, -0.3414264, -0.3414345, 
    -0.3413987, -0.3414252, -0.341428, -0.3414337, -0.3414352, -0.3414365, 
    -0.3414357, -0.3414315, -0.3414309, -0.341428, -0.3414271, -0.341425, 
    -0.3413976, -0.3414248, -0.3414265, -0.3414316, -0.341436, -0.341441, 
    -0.3414422, -0.3414477, -0.3414431, -0.3414505, -0.3414439, -0.3414554, 
    -0.3414352, -0.341444, -0.3414282, -0.3414299, -0.3414329, -0.3414401, 
    -0.3414364, -0.3414408, -0.3414308, -0.3414256, -0.3413987, -0.3413963, 
    -0.3413988, -0.3413986, -0.3414266, -0.3414259, -0.3414317, -0.3414286, 
    -0.3414375, -0.3414408, -0.34145, -0.3414556, -0.3414615, -0.341464, 
    -0.3414648, -0.3414652 ;

 TAUY =
  -0.341361, -0.3413828, -0.3413818, -0.3413859, -0.3413837, -0.3413863, 
    -0.3413621, -0.3413829, -0.3413637, -0.3413616, -0.3413936, -0.3413861, 
    -0.3414276, -0.341397, -0.3414353, -0.3414268, -0.3414371, -0.3414352, 
    -0.3414412, -0.3414395, -0.3414468, -0.3414419, -0.3414508, -0.3414457, 
    -0.3414465, -0.3414418, -0.3413877, -0.3413927, -0.3413874, -0.3413881, 
    -0.3413878, -0.3413837, -0.3413815, -0.3413607, -0.3413615, -0.3413812, 
    -0.3413884, -0.341386, -0.3413922, -0.3413921, -0.3413989, -0.3413958, 
    -0.3414331, -0.3414298, -0.3414395, -0.3414371, -0.3414394, -0.3414387, 
    -0.3414394, -0.3414358, -0.3414373, -0.3414342, -0.3413964, -0.3414255, 
    -0.3413894, -0.3413829, -0.3413623, -0.3413594, -0.3413598, -0.3413605, 
    -0.3413812, -0.3413852, -0.3413882, -0.3413901, -0.3413921, -0.3413977, 
    -0.3414266, -0.3414338, -0.3414326, -0.3414347, -0.3414368, -0.3414403, 
    -0.3414398, -0.3414413, -0.3414347, -0.341439, -0.3414319, -0.3414338, 
    -0.3413922, -0.3413867, -0.341384, -0.341382, -0.3413601, -0.3413637, 
    -0.3413623, -0.3413824, -0.3413846, -0.3413835, -0.3413902, -0.3413876, 
    -0.3414268, -0.3413953, -0.3414366, -0.3414328, -0.3414375, -0.3414351, 
    -0.3414392, -0.3414355, -0.3414419, -0.3414432, -0.3414423, -0.341446, 
    -0.3414353, -0.3414394, -0.3413835, -0.3413836, -0.3413845, -0.3413807, 
    -0.341364, -0.3413607, -0.3413636, -0.3413815, -0.3413847, -0.3413866, 
    -0.3413883, -0.3413923, -0.3413966, -0.3414285, -0.341433, -0.3414361, 
    -0.3414343, -0.3414359, -0.3414341, -0.3414332, -0.3414427, -0.3414373, 
    -0.3414454, -0.341445, -0.3414413, -0.341445, -0.3413838, -0.3413827, 
    -0.3413626, -0.341382, -0.3413603, -0.3413631, -0.3413813, -0.3413875, 
    -0.341389, -0.3413903, -0.3413928, -0.341396, -0.3414272, -0.3414323, 
    -0.341437, -0.3414367, -0.3414367, -0.3414378, -0.3414352, -0.3414382, 
    -0.3414387, -0.3414374, -0.3414449, -0.3414428, -0.341445, -0.3414436, 
    -0.3413831, -0.3413848, -0.3413838, -0.3413856, -0.3413843, -0.3413897, 
    -0.3413913, -0.3413989, -0.3413959, -0.3414265, -0.3413964, -0.3413972, 
    -0.3414265, -0.3413967, -0.3414319, -0.3414252, -0.3414378, -0.3414309, 
    -0.3414382, -0.341437, -0.3414391, -0.3414409, -0.3414434, -0.3414477, 
    -0.3414467, -0.3414504, -0.3413873, -0.3413895, -0.3413894, -0.3413917, 
    -0.3413934, -0.3413971, -0.3414287, -0.3414265, -0.3414307, -0.3414315, 
    -0.3414251, -0.341429, -0.341391, -0.3413929, -0.3413918, -0.3413875, 
    -0.3414269, -0.3413941, -0.3414331, -0.3414292, -0.3414407, -0.3414349, 
    -0.3414462, -0.3414508, -0.3414555, -0.3414606, -0.3413907, -0.3413893, 
    -0.341392, -0.3413956, -0.3414247, -0.3414294, -0.3414299, -0.3414308, 
    -0.3414331, -0.341435, -0.341431, -0.3414355, -0.3413932, -0.3414275, 
    -0.3413886, -0.3413925, -0.3413954, -0.3413942, -0.3414262, -0.3414277, 
    -0.3414339, -0.3414307, -0.3414496, -0.3414412, -0.3414647, -0.3414581, 
    -0.3413887, -0.3413908, -0.3413977, -0.3413944, -0.3414298, -0.3414322, 
    -0.3414342, -0.3414366, -0.341437, -0.3414384, -0.341436, -0.3414383, 
    -0.3414294, -0.3414334, -0.341397, -0.3414252, -0.3413984, -0.3413971, 
    -0.3414268, -0.3414311, -0.3414313, -0.3414326, -0.3414362, -0.3414298, 
    -0.3414505, -0.3414375, -0.341393, -0.3413967, -0.3413974, -0.3413959, 
    -0.3414319, -0.3414281, -0.3414384, -0.3414356, -0.3414402, -0.3414379, 
    -0.3414376, -0.3414347, -0.3414329, -0.3414283, -0.341399, -0.3413962, 
    -0.3413968, -0.3414255, -0.3414313, -0.3414369, -0.3414357, -0.3414398, 
    -0.3414291, -0.3414335, -0.3414317, -0.3414364, -0.3414264, -0.3414345, 
    -0.3413987, -0.3414252, -0.341428, -0.3414337, -0.3414352, -0.3414365, 
    -0.3414357, -0.3414315, -0.3414309, -0.341428, -0.3414271, -0.341425, 
    -0.3413976, -0.3414248, -0.3414265, -0.3414316, -0.341436, -0.341441, 
    -0.3414422, -0.3414477, -0.3414431, -0.3414505, -0.3414439, -0.3414554, 
    -0.3414352, -0.341444, -0.3414282, -0.3414299, -0.3414329, -0.3414401, 
    -0.3414364, -0.3414408, -0.3414308, -0.3414256, -0.3413987, -0.3413963, 
    -0.3413988, -0.3413986, -0.3414266, -0.3414259, -0.3414317, -0.3414286, 
    -0.3414375, -0.3414408, -0.34145, -0.3414556, -0.3414615, -0.341464, 
    -0.3414648, -0.3414652 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.7202, 261.7405, 261.7365, 261.753, 261.7439, 261.7547, 261.7243, 
    261.7413, 261.7305, 261.722, 261.7849, 261.7538, 261.8169, 261.7975, 
    261.847, 261.8138, 261.8537, 261.846, 261.869, 261.8624, 261.8918, 
    261.872, 261.907, 261.8871, 261.8902, 261.8714, 261.76, 261.781, 
    261.7588, 261.7618, 261.7604, 261.7441, 261.7358, 261.7186, 261.7217, 
    261.7343, 261.7631, 261.7534, 261.778, 261.7774, 261.8048, 261.7925, 
    261.838, 261.825, 261.8627, 261.8532, 261.8622, 261.8595, 261.8623, 
    261.8484, 261.8543, 261.8421, 261.7948, 261.8084, 261.7669, 261.7417, 
    261.725, 261.7132, 261.7148, 261.718, 261.7344, 261.7499, 261.7617, 
    261.7696, 261.7773, 261.8008, 261.8128, 261.8407, 261.8357, 261.8441, 
    261.8523, 261.8659, 261.8636, 261.8697, 261.8439, 261.861, 261.8328, 
    261.8405, 261.7794, 261.756, 261.746, 261.7373, 261.7161, 261.7308, 
    261.725, 261.7387, 261.7475, 261.7431, 261.7698, 261.7594, 261.8136, 
    261.7905, 261.8513, 261.8367, 261.8548, 261.8456, 261.8614, 261.8472, 
    261.8719, 261.8773, 261.8736, 261.8877, 261.8464, 261.8622, 261.743, 
    261.7437, 261.747, 261.7325, 261.7318, 261.7185, 261.7303, 261.7352, 
    261.748, 261.7555, 261.7626, 261.7784, 261.7959, 261.82, 261.8376, 
    261.8494, 261.8422, 261.8486, 261.8415, 261.8381, 261.8752, 261.8544, 
    261.8857, 261.884, 261.8698, 261.8842, 261.7442, 261.7401, 261.7261, 
    261.7371, 261.7171, 261.7283, 261.7347, 261.7596, 261.7651, 261.7702, 
    261.7802, 261.7931, 261.8152, 261.8348, 261.8528, 261.8514, 261.8519, 
    261.8559, 261.846, 261.8575, 261.8594, 261.8544, 261.8837, 261.8753, 
    261.8839, 261.8785, 261.7415, 261.7483, 261.7446, 261.7516, 261.7466, 
    261.7684, 261.7749, 261.8053, 261.7928, 261.8123, 261.7949, 261.798, 
    261.8129, 261.7958, 261.8337, 261.8077, 261.856, 261.8301, 261.8577, 
    261.8527, 261.861, 261.8684, 261.8777, 261.8949, 261.8909, 261.9053, 
    261.7585, 261.7673, 261.7665, 261.7758, 261.7827, 261.7975, 261.8208, 
    261.8119, 261.8283, 261.8316, 261.8067, 261.822, 261.7733, 261.7812, 
    261.7765, 261.7592, 261.8139, 261.786, 261.8379, 261.8226, 261.8673, 
    261.8451, 261.8887, 261.9073, 261.9249, 261.9454, 261.7722, 261.7661, 
    261.7769, 261.7918, 261.8052, 261.8235, 261.8254, 261.8288, 261.8377, 
    261.8452, 261.8299, 261.8471, 261.783, 261.8164, 261.7639, 261.7798, 
    261.7909, 261.786, 261.8109, 261.8168, 261.841, 261.8285, 261.9027, 
    261.8699, 261.961, 261.9355, 261.764, 261.7721, 261.8003, 261.7869, 
    261.8248, 261.8342, 261.8418, 261.8516, 261.8527, 261.8585, 261.849, 
    261.8581, 261.8236, 261.839, 261.7971, 261.8069, 261.8026, 261.7974, 
    261.8131, 261.8301, 261.8305, 261.836, 261.8514, 261.8249, 261.907, 
    261.8563, 261.7809, 261.7965, 261.7988, 261.7927, 261.8332, 261.8184, 
    261.8583, 261.8475, 261.8652, 261.8564, 261.8551, 261.8438, 261.8368, 
    261.8191, 261.8051, 261.7936, 261.7963, 261.8084, 261.8312, 261.8528, 
    261.848, 261.8639, 261.822, 261.8395, 261.8327, 261.8505, 261.8117, 
    261.8446, 261.8036, 261.8069, 261.8181, 261.8407, 261.8457, 261.8511, 
    261.8478, 261.8318, 261.8292, 261.8178, 261.8147, 261.8061, 261.7993, 
    261.8055, 261.8123, 261.8318, 261.8493, 261.8685, 261.8732, 261.8954, 
    261.8773, 261.9072, 261.8817, 261.9259, 261.8466, 261.881, 261.8186, 
    261.8253, 261.8375, 261.8654, 261.8504, 261.868, 261.8291, 261.8088, 
    261.804, 261.7943, 261.8043, 261.8035, 261.8126, 261.8095, 261.8325, 
    261.8201, 261.8551, 261.8678, 261.9038, 261.9258, 261.9482, 261.9581, 
    261.9612, 261.9624 ;

 TG_R =
  261.7202, 261.7405, 261.7365, 261.753, 261.7439, 261.7547, 261.7243, 
    261.7413, 261.7305, 261.722, 261.7849, 261.7538, 261.8169, 261.7975, 
    261.847, 261.8138, 261.8537, 261.846, 261.869, 261.8624, 261.8918, 
    261.872, 261.907, 261.8871, 261.8902, 261.8714, 261.76, 261.781, 
    261.7588, 261.7618, 261.7604, 261.7441, 261.7358, 261.7186, 261.7217, 
    261.7343, 261.7631, 261.7534, 261.778, 261.7774, 261.8048, 261.7925, 
    261.838, 261.825, 261.8627, 261.8532, 261.8622, 261.8595, 261.8623, 
    261.8484, 261.8543, 261.8421, 261.7948, 261.8084, 261.7669, 261.7417, 
    261.725, 261.7132, 261.7148, 261.718, 261.7344, 261.7499, 261.7617, 
    261.7696, 261.7773, 261.8008, 261.8128, 261.8407, 261.8357, 261.8441, 
    261.8523, 261.8659, 261.8636, 261.8697, 261.8439, 261.861, 261.8328, 
    261.8405, 261.7794, 261.756, 261.746, 261.7373, 261.7161, 261.7308, 
    261.725, 261.7387, 261.7475, 261.7431, 261.7698, 261.7594, 261.8136, 
    261.7905, 261.8513, 261.8367, 261.8548, 261.8456, 261.8614, 261.8472, 
    261.8719, 261.8773, 261.8736, 261.8877, 261.8464, 261.8622, 261.743, 
    261.7437, 261.747, 261.7325, 261.7318, 261.7185, 261.7303, 261.7352, 
    261.748, 261.7555, 261.7626, 261.7784, 261.7959, 261.82, 261.8376, 
    261.8494, 261.8422, 261.8486, 261.8415, 261.8381, 261.8752, 261.8544, 
    261.8857, 261.884, 261.8698, 261.8842, 261.7442, 261.7401, 261.7261, 
    261.7371, 261.7171, 261.7283, 261.7347, 261.7596, 261.7651, 261.7702, 
    261.7802, 261.7931, 261.8152, 261.8348, 261.8528, 261.8514, 261.8519, 
    261.8559, 261.846, 261.8575, 261.8594, 261.8544, 261.8837, 261.8753, 
    261.8839, 261.8785, 261.7415, 261.7483, 261.7446, 261.7516, 261.7466, 
    261.7684, 261.7749, 261.8053, 261.7928, 261.8123, 261.7949, 261.798, 
    261.8129, 261.7958, 261.8337, 261.8077, 261.856, 261.8301, 261.8577, 
    261.8527, 261.861, 261.8684, 261.8777, 261.8949, 261.8909, 261.9053, 
    261.7585, 261.7673, 261.7665, 261.7758, 261.7827, 261.7975, 261.8208, 
    261.8119, 261.8283, 261.8316, 261.8067, 261.822, 261.7733, 261.7812, 
    261.7765, 261.7592, 261.8139, 261.786, 261.8379, 261.8226, 261.8673, 
    261.8451, 261.8887, 261.9073, 261.9249, 261.9454, 261.7722, 261.7661, 
    261.7769, 261.7918, 261.8052, 261.8235, 261.8254, 261.8288, 261.8377, 
    261.8452, 261.8299, 261.8471, 261.783, 261.8164, 261.7639, 261.7798, 
    261.7909, 261.786, 261.8109, 261.8168, 261.841, 261.8285, 261.9027, 
    261.8699, 261.961, 261.9355, 261.764, 261.7721, 261.8003, 261.7869, 
    261.8248, 261.8342, 261.8418, 261.8516, 261.8527, 261.8585, 261.849, 
    261.8581, 261.8236, 261.839, 261.7971, 261.8069, 261.8026, 261.7974, 
    261.8131, 261.8301, 261.8305, 261.836, 261.8514, 261.8249, 261.907, 
    261.8563, 261.7809, 261.7965, 261.7988, 261.7927, 261.8332, 261.8184, 
    261.8583, 261.8475, 261.8652, 261.8564, 261.8551, 261.8438, 261.8368, 
    261.8191, 261.8051, 261.7936, 261.7963, 261.8084, 261.8312, 261.8528, 
    261.848, 261.8639, 261.822, 261.8395, 261.8327, 261.8505, 261.8117, 
    261.8446, 261.8036, 261.8069, 261.8181, 261.8407, 261.8457, 261.8511, 
    261.8478, 261.8318, 261.8292, 261.8178, 261.8147, 261.8061, 261.7993, 
    261.8055, 261.8123, 261.8318, 261.8493, 261.8685, 261.8732, 261.8954, 
    261.8773, 261.9072, 261.8817, 261.9259, 261.8466, 261.881, 261.8186, 
    261.8253, 261.8375, 261.8654, 261.8504, 261.868, 261.8291, 261.8088, 
    261.804, 261.7943, 261.8043, 261.8035, 261.8126, 261.8095, 261.8325, 
    261.8201, 261.8551, 261.8678, 261.9038, 261.9258, 261.9482, 261.9581, 
    261.9612, 261.9624 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.6766, 254.6781, 254.6778, 254.6791, 254.6784, 254.6792, 254.6769, 
    254.6782, 254.6774, 254.6768, 254.6814, 254.6791, 254.6839, 254.6824, 
    254.6862, 254.6837, 254.6867, 254.6861, 254.6879, 254.6874, 254.6896, 
    254.6881, 254.6908, 254.6893, 254.6895, 254.6881, 254.6796, 254.6811, 
    254.6795, 254.6797, 254.6796, 254.6784, 254.6778, 254.6765, 254.6767, 
    254.6777, 254.6798, 254.6791, 254.681, 254.6809, 254.683, 254.6821, 
    254.6855, 254.6846, 254.6874, 254.6867, 254.6874, 254.6872, 254.6874, 
    254.6863, 254.6868, 254.6858, 254.6822, 254.6833, 254.6801, 254.6782, 
    254.677, 254.6761, 254.6762, 254.6765, 254.6777, 254.6788, 254.6797, 
    254.6803, 254.6809, 254.6826, 254.6836, 254.6857, 254.6854, 254.686, 
    254.6866, 254.6877, 254.6875, 254.6879, 254.686, 254.6873, 254.6852, 
    254.6857, 254.681, 254.6793, 254.6785, 254.6779, 254.6763, 254.6774, 
    254.677, 254.678, 254.6787, 254.6783, 254.6803, 254.6796, 254.6837, 
    254.6819, 254.6865, 254.6854, 254.6868, 254.6861, 254.6873, 254.6862, 
    254.6881, 254.6885, 254.6882, 254.6893, 254.6862, 254.6874, 254.6783, 
    254.6784, 254.6786, 254.6775, 254.6775, 254.6765, 254.6774, 254.6777, 
    254.6787, 254.6793, 254.6798, 254.681, 254.6823, 254.6842, 254.6855, 
    254.6864, 254.6859, 254.6863, 254.6858, 254.6855, 254.6884, 254.6868, 
    254.6892, 254.689, 254.6879, 254.689, 254.6784, 254.6781, 254.6771, 
    254.6779, 254.6764, 254.6772, 254.6777, 254.6796, 254.68, 254.6804, 
    254.6811, 254.6821, 254.6838, 254.6853, 254.6867, 254.6866, 254.6866, 
    254.6869, 254.6861, 254.687, 254.6871, 254.6868, 254.689, 254.6884, 
    254.689, 254.6886, 254.6782, 254.6787, 254.6785, 254.679, 254.6786, 
    254.6802, 254.6807, 254.683, 254.6821, 254.6836, 254.6822, 254.6825, 
    254.6836, 254.6823, 254.6852, 254.6832, 254.6869, 254.6849, 254.687, 
    254.6866, 254.6873, 254.6878, 254.6886, 254.6898, 254.6896, 254.6907, 
    254.6795, 254.6801, 254.6801, 254.6808, 254.6813, 254.6824, 254.6842, 
    254.6836, 254.6848, 254.685, 254.6832, 254.6843, 254.6806, 254.6812, 
    254.6808, 254.6795, 254.6837, 254.6815, 254.6855, 254.6844, 254.6878, 
    254.6861, 254.6894, 254.6908, 254.6922, 254.6937, 254.6805, 254.6801, 
    254.6809, 254.682, 254.683, 254.6844, 254.6846, 254.6848, 254.6855, 
    254.6861, 254.6849, 254.6862, 254.6813, 254.6839, 254.6799, 254.6811, 
    254.6819, 254.6816, 254.6835, 254.6839, 254.6857, 254.6848, 254.6904, 
    254.6879, 254.6949, 254.6929, 254.6799, 254.6805, 254.6826, 254.6816, 
    254.6845, 254.6852, 254.6858, 254.6866, 254.6866, 254.6871, 254.6864, 
    254.6871, 254.6844, 254.6856, 254.6824, 254.6832, 254.6828, 254.6824, 
    254.6837, 254.6849, 254.685, 254.6854, 254.6865, 254.6845, 254.6907, 
    254.6869, 254.6812, 254.6823, 254.6825, 254.6821, 254.6852, 254.6841, 
    254.6871, 254.6863, 254.6876, 254.6869, 254.6868, 254.686, 254.6854, 
    254.6841, 254.683, 254.6821, 254.6823, 254.6833, 254.685, 254.6866, 
    254.6863, 254.6875, 254.6843, 254.6856, 254.6851, 254.6865, 254.6835, 
    254.686, 254.6829, 254.6832, 254.684, 254.6857, 254.6861, 254.6865, 
    254.6863, 254.6851, 254.6849, 254.684, 254.6838, 254.6831, 254.6826, 
    254.6831, 254.6836, 254.6851, 254.6864, 254.6878, 254.6882, 254.6899, 
    254.6885, 254.6907, 254.6888, 254.6922, 254.6862, 254.6888, 254.6841, 
    254.6846, 254.6855, 254.6876, 254.6865, 254.6878, 254.6849, 254.6833, 
    254.6829, 254.6822, 254.683, 254.6829, 254.6836, 254.6834, 254.6851, 
    254.6842, 254.6868, 254.6878, 254.6905, 254.6922, 254.6939, 254.6947, 
    254.6949, 254.695 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.2395, 18.23949, 18.23949, 18.23948, 18.23949, 18.23948, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23947, 18.23948, 18.23945, 18.23946, 
    18.23944, 18.23945, 18.23944, 18.23944, 18.23943, 18.23943, 18.23942, 
    18.23943, 18.23941, 18.23942, 18.23942, 18.23943, 18.23948, 18.23947, 
    18.23948, 18.23948, 18.23948, 18.23949, 18.23949, 18.2395, 18.2395, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23947, 
    18.23944, 18.23945, 18.23943, 18.23944, 18.23943, 18.23943, 18.23943, 
    18.23944, 18.23944, 18.23944, 18.23946, 18.23946, 18.23948, 18.23949, 
    18.2395, 18.2395, 18.2395, 18.2395, 18.23949, 18.23949, 18.23948, 
    18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23943, 18.23943, 18.23943, 18.23944, 18.23943, 18.23944, 
    18.23944, 18.23947, 18.23948, 18.23949, 18.23949, 18.2395, 18.2395, 
    18.2395, 18.23949, 18.23949, 18.23949, 18.23948, 18.23948, 18.23945, 
    18.23947, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23942, 18.23943, 18.23942, 18.23944, 18.23943, 18.23949, 
    18.23949, 18.23949, 18.23949, 18.23949, 18.2395, 18.2395, 18.23949, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23944, 18.23944, 18.23944, 18.23944, 18.23942, 18.23944, 
    18.23942, 18.23942, 18.23943, 18.23942, 18.23949, 18.23949, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23949, 18.23948, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23942, 18.23942, 
    18.23942, 18.23942, 18.23949, 18.23949, 18.23949, 18.23948, 18.23949, 
    18.23948, 18.23947, 18.23946, 18.23947, 18.23946, 18.23946, 18.23946, 
    18.23945, 18.23946, 18.23944, 18.23946, 18.23943, 18.23945, 18.23943, 
    18.23944, 18.23943, 18.23943, 18.23942, 18.23941, 18.23942, 18.23941, 
    18.23948, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23945, 
    18.23946, 18.23945, 18.23945, 18.23946, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23948, 18.23945, 18.23947, 18.23944, 18.23945, 18.23943, 
    18.23944, 18.23942, 18.23941, 18.2394, 18.23939, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23945, 18.23945, 18.23944, 
    18.23944, 18.23945, 18.23944, 18.23947, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23938, 18.2394, 18.23948, 18.23948, 18.23946, 18.23947, 
    18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23945, 18.23944, 18.23946, 18.23946, 18.23946, 18.23946, 
    18.23945, 18.23945, 18.23945, 18.23944, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23947, 18.23946, 18.23946, 18.23947, 18.23944, 18.23945, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23944, 18.23944, 
    18.23945, 18.23946, 18.23947, 18.23946, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23943, 18.23945, 18.23944, 18.23944, 18.23944, 18.23946, 
    18.23944, 18.23946, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23945, 18.23945, 18.23945, 18.23945, 18.23946, 18.23946, 
    18.23946, 18.23946, 18.23945, 18.23944, 18.23943, 18.23943, 18.23941, 
    18.23942, 18.23941, 18.23942, 18.2394, 18.23944, 18.23942, 18.23945, 
    18.23945, 18.23944, 18.23943, 18.23944, 18.23943, 18.23945, 18.23946, 
    18.23946, 18.23946, 18.23946, 18.23946, 18.23946, 18.23946, 18.23944, 
    18.23945, 18.23944, 18.23943, 18.23941, 18.2394, 18.23939, 18.23938, 
    18.23938, 18.23938 ;

 TOTCOLCH4 =
  1.320645e-05, 1.302424e-05, 1.305964e-05, 1.291288e-05, 1.299427e-05, 
    1.289821e-05, 1.316949e-05, 1.3017e-05, 1.311432e-05, 1.319005e-05, 
    1.262882e-05, 1.290635e-05, 1.234172e-05, 1.251791e-05, 1.207616e-05, 
    1.236909e-05, 1.201725e-05, 1.208462e-05, 1.188213e-05, 1.194008e-05, 
    1.168171e-05, 1.18554e-05, 1.154823e-05, 1.172316e-05, 1.169575e-05, 
    1.186113e-05, 1.285044e-05, 1.266331e-05, 1.286154e-05, 1.283482e-05, 
    1.284681e-05, 1.299258e-05, 1.306611e-05, 1.322041e-05, 1.319238e-05, 
    1.307908e-05, 1.282281e-05, 1.290973e-05, 1.269091e-05, 1.269585e-05, 
    1.245294e-05, 1.256236e-05, 1.21553e-05, 1.227076e-05, 1.193766e-05, 
    1.202127e-05, 1.194158e-05, 1.196574e-05, 1.194126e-05, 1.206394e-05, 
    1.201135e-05, 1.21194e-05, 1.254185e-05, 1.241743e-05, 1.278911e-05, 
    1.301341e-05, 1.316279e-05, 1.326893e-05, 1.325392e-05, 1.32253e-05, 
    1.307841e-05, 1.294056e-05, 1.283566e-05, 1.276556e-05, 1.269656e-05, 
    1.2488e-05, 1.23779e-05, 1.213196e-05, 1.217631e-05, 1.210122e-05, 
    1.20296e-05, 1.190949e-05, 1.192925e-05, 1.187638e-05, 1.210322e-05, 
    1.195237e-05, 1.220157e-05, 1.213332e-05, 1.267772e-05, 1.288628e-05, 
    1.297501e-05, 1.305283e-05, 1.324238e-05, 1.311143e-05, 1.316302e-05, 
    1.304035e-05, 1.296248e-05, 1.300098e-05, 1.276365e-05, 1.285583e-05, 
    1.237138e-05, 1.257967e-05, 1.203795e-05, 1.21672e-05, 1.200701e-05, 
    1.208871e-05, 1.194877e-05, 1.20747e-05, 1.185672e-05, 1.180935e-05, 
    1.184172e-05, 1.171749e-05, 1.208169e-05, 1.194157e-05, 1.300206e-05, 
    1.299578e-05, 1.296652e-05, 1.309518e-05, 1.310306e-05, 1.322117e-05, 
    1.311608e-05, 1.307136e-05, 1.295797e-05, 1.289096e-05, 1.282732e-05, 
    1.268757e-05, 1.253177e-05, 1.23145e-05, 1.215882e-05, 1.205465e-05, 
    1.211851e-05, 1.206213e-05, 1.212516e-05, 1.215472e-05, 1.182709e-05, 
    1.201085e-05, 1.173534e-05, 1.175056e-05, 1.187512e-05, 1.174884e-05, 
    1.299137e-05, 1.302752e-05, 1.315314e-05, 1.305481e-05, 1.323405e-05, 
    1.313366e-05, 1.307599e-05, 1.285388e-05, 1.280519e-05, 1.276003e-05, 
    1.267095e-05, 1.255676e-05, 1.235686e-05, 1.21834e-05, 1.202544e-05, 
    1.2037e-05, 1.203293e-05, 1.199768e-05, 1.208502e-05, 1.198335e-05, 
    1.19663e-05, 1.201089e-05, 1.17526e-05, 1.182628e-05, 1.175088e-05, 
    1.179885e-05, 1.301577e-05, 1.295496e-05, 1.298781e-05, 1.292604e-05, 
    1.296955e-05, 1.277624e-05, 1.271838e-05, 1.244822e-05, 1.2559e-05, 
    1.23828e-05, 1.254109e-05, 1.251301e-05, 1.237702e-05, 1.253253e-05, 
    1.219293e-05, 1.242296e-05, 1.199631e-05, 1.222533e-05, 1.198198e-05, 
    1.202612e-05, 1.195306e-05, 1.188769e-05, 1.180557e-05, 1.165428e-05, 
    1.168928e-05, 1.156299e-05, 1.286439e-05, 1.278567e-05, 1.279261e-05, 
    1.271031e-05, 1.26495e-05, 1.251788e-05, 1.230724e-05, 1.238638e-05, 
    1.224118e-05, 1.221206e-05, 1.243269e-05, 1.229713e-05, 1.273303e-05, 
    1.266242e-05, 1.270447e-05, 1.285817e-05, 1.236811e-05, 1.261921e-05, 
    1.215624e-05, 1.229176e-05, 1.189701e-05, 1.209302e-05, 1.170856e-05, 
    1.154486e-05, 1.139128e-05, 1.121223e-05, 1.274275e-05, 1.27962e-05, 
    1.270053e-05, 1.256833e-05, 1.244593e-05, 1.228349e-05, 1.22669e-05, 
    1.223651e-05, 1.215787e-05, 1.209182e-05, 1.222689e-05, 1.207527e-05, 
    1.264602e-05, 1.234637e-05, 1.281641e-05, 1.267454e-05, 1.257613e-05, 
    1.26193e-05, 1.239544e-05, 1.234277e-05, 1.212914e-05, 1.22395e-05, 
    1.158521e-05, 1.187387e-05, 1.107632e-05, 1.129811e-05, 1.281489e-05, 
    1.274294e-05, 1.249305e-05, 1.261185e-05, 1.227266e-05, 1.218941e-05, 
    1.212182e-05, 1.203549e-05, 1.202619e-05, 1.19751e-05, 1.205884e-05, 
    1.197841e-05, 1.228314e-05, 1.21468e-05, 1.252159e-05, 1.243018e-05, 
    1.247223e-05, 1.251836e-05, 1.237607e-05, 1.222475e-05, 1.222155e-05, 
    1.21731e-05, 1.20367e-05, 1.227129e-05, 1.1548e-05, 1.19937e-05, 
    1.266457e-05, 1.252629e-05, 1.250659e-05, 1.25601e-05, 1.219775e-05, 
    1.232883e-05, 1.197635e-05, 1.207144e-05, 1.191571e-05, 1.199305e-05, 
    1.200443e-05, 1.210391e-05, 1.216591e-05, 1.232281e-05, 1.245073e-05, 
    1.255234e-05, 1.252871e-05, 1.241713e-05, 1.221551e-05, 1.202533e-05, 
    1.206694e-05, 1.192753e-05, 1.22972e-05, 1.214194e-05, 1.22019e-05, 
    1.204567e-05, 1.238848e-05, 1.209637e-05, 1.246333e-05, 1.243109e-05, 
    1.233144e-05, 1.21314e-05, 1.208726e-05, 1.204012e-05, 1.206921e-05, 
    1.221041e-05, 1.223358e-05, 1.233386e-05, 1.236156e-05, 1.243811e-05, 
    1.250153e-05, 1.244357e-05, 1.238276e-05, 1.221036e-05, 1.205535e-05, 
    1.188676e-05, 1.184558e-05, 1.164922e-05, 1.180898e-05, 1.154552e-05, 
    1.176939e-05, 1.138241e-05, 1.207952e-05, 1.177604e-05, 1.232691e-05, 
    1.226736e-05, 1.215974e-05, 1.191361e-05, 1.20464e-05, 1.189114e-05, 
    1.223449e-05, 1.241327e-05, 1.245963e-05, 1.254616e-05, 1.245766e-05, 
    1.246485e-05, 1.238026e-05, 1.240743e-05, 1.220464e-05, 1.23135e-05, 
    1.200471e-05, 1.189237e-05, 1.15762e-05, 1.138317e-05, 1.118736e-05, 
    1.110112e-05, 1.10749e-05, 1.106394e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.2395, 18.23949, 18.23949, 18.23948, 18.23949, 18.23948, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23947, 18.23948, 18.23945, 18.23946, 
    18.23944, 18.23945, 18.23944, 18.23944, 18.23943, 18.23943, 18.23942, 
    18.23943, 18.23941, 18.23942, 18.23942, 18.23943, 18.23948, 18.23947, 
    18.23948, 18.23948, 18.23948, 18.23949, 18.23949, 18.2395, 18.2395, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23947, 
    18.23944, 18.23945, 18.23943, 18.23944, 18.23943, 18.23943, 18.23943, 
    18.23944, 18.23944, 18.23944, 18.23946, 18.23946, 18.23948, 18.23949, 
    18.2395, 18.2395, 18.2395, 18.2395, 18.23949, 18.23949, 18.23948, 
    18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23943, 18.23943, 18.23943, 18.23944, 18.23943, 18.23944, 
    18.23944, 18.23947, 18.23948, 18.23949, 18.23949, 18.2395, 18.2395, 
    18.2395, 18.23949, 18.23949, 18.23949, 18.23948, 18.23948, 18.23945, 
    18.23947, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23942, 18.23943, 18.23942, 18.23944, 18.23943, 18.23949, 
    18.23949, 18.23949, 18.23949, 18.23949, 18.2395, 18.2395, 18.23949, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23944, 18.23944, 18.23944, 18.23944, 18.23942, 18.23944, 
    18.23942, 18.23942, 18.23943, 18.23942, 18.23949, 18.23949, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23949, 18.23948, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23942, 18.23942, 
    18.23942, 18.23942, 18.23949, 18.23949, 18.23949, 18.23948, 18.23949, 
    18.23948, 18.23947, 18.23946, 18.23947, 18.23946, 18.23946, 18.23946, 
    18.23945, 18.23946, 18.23944, 18.23946, 18.23943, 18.23945, 18.23943, 
    18.23944, 18.23943, 18.23943, 18.23942, 18.23941, 18.23942, 18.23941, 
    18.23948, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23945, 
    18.23946, 18.23945, 18.23945, 18.23946, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23948, 18.23945, 18.23947, 18.23944, 18.23945, 18.23943, 
    18.23944, 18.23942, 18.23941, 18.2394, 18.23939, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23945, 18.23945, 18.23944, 
    18.23944, 18.23945, 18.23944, 18.23947, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23938, 18.2394, 18.23948, 18.23948, 18.23946, 18.23947, 
    18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23945, 18.23944, 18.23946, 18.23946, 18.23946, 18.23946, 
    18.23945, 18.23945, 18.23945, 18.23944, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23947, 18.23946, 18.23946, 18.23947, 18.23944, 18.23945, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23944, 18.23944, 
    18.23945, 18.23946, 18.23947, 18.23946, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23943, 18.23945, 18.23944, 18.23944, 18.23944, 18.23946, 
    18.23944, 18.23946, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23945, 18.23945, 18.23945, 18.23945, 18.23946, 18.23946, 
    18.23946, 18.23946, 18.23945, 18.23944, 18.23943, 18.23943, 18.23941, 
    18.23942, 18.23941, 18.23942, 18.2394, 18.23944, 18.23942, 18.23945, 
    18.23945, 18.23944, 18.23943, 18.23944, 18.23943, 18.23945, 18.23946, 
    18.23946, 18.23946, 18.23946, 18.23946, 18.23946, 18.23946, 18.23944, 
    18.23945, 18.23944, 18.23943, 18.23941, 18.2394, 18.23939, 18.23938, 
    18.23938, 18.23938 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976081e-05, 5.976067e-05, 5.97607e-05, 5.976058e-05, 5.976064e-05, 
    5.976057e-05, 5.976078e-05, 5.976066e-05, 5.976074e-05, 5.97608e-05, 
    5.976036e-05, 5.976058e-05, 5.976013e-05, 5.976027e-05, 5.975992e-05, 
    5.976015e-05, 5.975987e-05, 5.975993e-05, 5.975977e-05, 5.975981e-05, 
    5.975961e-05, 5.975975e-05, 5.97595e-05, 5.975964e-05, 5.975962e-05, 
    5.975975e-05, 5.976053e-05, 5.976039e-05, 5.976054e-05, 5.976052e-05, 
    5.976053e-05, 5.976064e-05, 5.97607e-05, 5.976082e-05, 5.97608e-05, 
    5.976071e-05, 5.976051e-05, 5.976058e-05, 5.97604e-05, 5.976041e-05, 
    5.976022e-05, 5.976031e-05, 5.975998e-05, 5.976007e-05, 5.975981e-05, 
    5.975988e-05, 5.975981e-05, 5.975983e-05, 5.975981e-05, 5.975991e-05, 
    5.975987e-05, 5.975995e-05, 5.976029e-05, 5.976019e-05, 5.976048e-05, 
    5.976066e-05, 5.976078e-05, 5.976086e-05, 5.976085e-05, 5.976083e-05, 
    5.976071e-05, 5.97606e-05, 5.976052e-05, 5.976047e-05, 5.976041e-05, 
    5.976024e-05, 5.976016e-05, 5.975996e-05, 5.976e-05, 5.975994e-05, 
    5.975988e-05, 5.975979e-05, 5.97598e-05, 5.975976e-05, 5.975994e-05, 
    5.975982e-05, 5.976002e-05, 5.975996e-05, 5.97604e-05, 5.976056e-05, 
    5.976063e-05, 5.976069e-05, 5.976084e-05, 5.976074e-05, 5.976078e-05, 
    5.976068e-05, 5.976062e-05, 5.976065e-05, 5.976046e-05, 5.976054e-05, 
    5.976015e-05, 5.976032e-05, 5.975989e-05, 5.975999e-05, 5.975987e-05, 
    5.975993e-05, 5.975982e-05, 5.975992e-05, 5.975975e-05, 5.975971e-05, 
    5.975974e-05, 5.975964e-05, 5.975992e-05, 5.975981e-05, 5.976065e-05, 
    5.976065e-05, 5.976062e-05, 5.976072e-05, 5.976073e-05, 5.976082e-05, 
    5.976074e-05, 5.976071e-05, 5.976062e-05, 5.976056e-05, 5.976051e-05, 
    5.97604e-05, 5.976028e-05, 5.976011e-05, 5.975999e-05, 5.97599e-05, 
    5.975995e-05, 5.975991e-05, 5.975996e-05, 5.975998e-05, 5.975972e-05, 
    5.975987e-05, 5.975965e-05, 5.975966e-05, 5.975976e-05, 5.975966e-05, 
    5.976064e-05, 5.976067e-05, 5.976077e-05, 5.976069e-05, 5.976083e-05, 
    5.976075e-05, 5.976071e-05, 5.976054e-05, 5.97605e-05, 5.976046e-05, 
    5.976039e-05, 5.97603e-05, 5.976014e-05, 5.976e-05, 5.975988e-05, 
    5.975989e-05, 5.975988e-05, 5.975986e-05, 5.975993e-05, 5.975985e-05, 
    5.975983e-05, 5.975987e-05, 5.975966e-05, 5.975972e-05, 5.975966e-05, 
    5.97597e-05, 5.976066e-05, 5.976062e-05, 5.976064e-05, 5.976059e-05, 
    5.976063e-05, 5.976047e-05, 5.976043e-05, 5.976022e-05, 5.97603e-05, 
    5.976016e-05, 5.976029e-05, 5.976027e-05, 5.976016e-05, 5.976028e-05, 
    5.976001e-05, 5.976019e-05, 5.975986e-05, 5.976004e-05, 5.975984e-05, 
    5.975988e-05, 5.975982e-05, 5.975977e-05, 5.975971e-05, 5.975959e-05, 
    5.975961e-05, 5.975951e-05, 5.976054e-05, 5.976048e-05, 5.976049e-05, 
    5.976042e-05, 5.976037e-05, 5.976027e-05, 5.97601e-05, 5.976016e-05, 
    5.976005e-05, 5.976003e-05, 5.97602e-05, 5.97601e-05, 5.976044e-05, 
    5.976038e-05, 5.976042e-05, 5.976054e-05, 5.976015e-05, 5.976035e-05, 
    5.975998e-05, 5.976009e-05, 5.975978e-05, 5.975994e-05, 5.975963e-05, 
    5.97595e-05, 5.975938e-05, 5.975923e-05, 5.976045e-05, 5.976049e-05, 
    5.976042e-05, 5.976031e-05, 5.976021e-05, 5.976008e-05, 5.976007e-05, 
    5.976005e-05, 5.975999e-05, 5.975993e-05, 5.976004e-05, 5.975992e-05, 
    5.976037e-05, 5.976014e-05, 5.976051e-05, 5.976039e-05, 5.976032e-05, 
    5.976035e-05, 5.976017e-05, 5.976013e-05, 5.975996e-05, 5.976005e-05, 
    5.975953e-05, 5.975976e-05, 5.975912e-05, 5.97593e-05, 5.97605e-05, 
    5.976045e-05, 5.976025e-05, 5.976034e-05, 5.976008e-05, 5.976001e-05, 
    5.975996e-05, 5.975989e-05, 5.975988e-05, 5.975984e-05, 5.975991e-05, 
    5.975984e-05, 5.976008e-05, 5.975998e-05, 5.976027e-05, 5.97602e-05, 
    5.976023e-05, 5.976027e-05, 5.976016e-05, 5.976004e-05, 5.976003e-05, 
    5.976e-05, 5.975989e-05, 5.976007e-05, 5.97595e-05, 5.975986e-05, 
    5.976039e-05, 5.976028e-05, 5.976026e-05, 5.97603e-05, 5.976002e-05, 
    5.976012e-05, 5.975984e-05, 5.975992e-05, 5.975979e-05, 5.975986e-05, 
    5.975986e-05, 5.975994e-05, 5.975999e-05, 5.976012e-05, 5.976022e-05, 
    5.97603e-05, 5.976028e-05, 5.976019e-05, 5.976003e-05, 5.975988e-05, 
    5.975991e-05, 5.97598e-05, 5.97601e-05, 5.975997e-05, 5.976002e-05, 
    5.97599e-05, 5.976017e-05, 5.975994e-05, 5.976023e-05, 5.97602e-05, 
    5.976012e-05, 5.975996e-05, 5.975993e-05, 5.975989e-05, 5.975991e-05, 
    5.976003e-05, 5.976004e-05, 5.976012e-05, 5.976015e-05, 5.976021e-05, 
    5.976026e-05, 5.976021e-05, 5.976016e-05, 5.976003e-05, 5.97599e-05, 
    5.975977e-05, 5.975974e-05, 5.975958e-05, 5.975971e-05, 5.97595e-05, 
    5.975968e-05, 5.975937e-05, 5.975992e-05, 5.975968e-05, 5.976012e-05, 
    5.976007e-05, 5.975999e-05, 5.975979e-05, 5.97599e-05, 5.975978e-05, 
    5.976004e-05, 5.976019e-05, 5.976022e-05, 5.976029e-05, 5.976022e-05, 
    5.976023e-05, 5.976016e-05, 5.976018e-05, 5.976002e-05, 5.976011e-05, 
    5.975986e-05, 5.975978e-05, 5.975952e-05, 5.975937e-05, 5.975921e-05, 
    5.975914e-05, 5.975912e-05, 5.975911e-05 ;

 TOTLITC_1m =
  5.976081e-05, 5.976067e-05, 5.97607e-05, 5.976058e-05, 5.976064e-05, 
    5.976057e-05, 5.976078e-05, 5.976066e-05, 5.976074e-05, 5.97608e-05, 
    5.976036e-05, 5.976058e-05, 5.976013e-05, 5.976027e-05, 5.975992e-05, 
    5.976015e-05, 5.975987e-05, 5.975993e-05, 5.975977e-05, 5.975981e-05, 
    5.975961e-05, 5.975975e-05, 5.97595e-05, 5.975964e-05, 5.975962e-05, 
    5.975975e-05, 5.976053e-05, 5.976039e-05, 5.976054e-05, 5.976052e-05, 
    5.976053e-05, 5.976064e-05, 5.97607e-05, 5.976082e-05, 5.97608e-05, 
    5.976071e-05, 5.976051e-05, 5.976058e-05, 5.97604e-05, 5.976041e-05, 
    5.976022e-05, 5.976031e-05, 5.975998e-05, 5.976007e-05, 5.975981e-05, 
    5.975988e-05, 5.975981e-05, 5.975983e-05, 5.975981e-05, 5.975991e-05, 
    5.975987e-05, 5.975995e-05, 5.976029e-05, 5.976019e-05, 5.976048e-05, 
    5.976066e-05, 5.976078e-05, 5.976086e-05, 5.976085e-05, 5.976083e-05, 
    5.976071e-05, 5.97606e-05, 5.976052e-05, 5.976047e-05, 5.976041e-05, 
    5.976024e-05, 5.976016e-05, 5.975996e-05, 5.976e-05, 5.975994e-05, 
    5.975988e-05, 5.975979e-05, 5.97598e-05, 5.975976e-05, 5.975994e-05, 
    5.975982e-05, 5.976002e-05, 5.975996e-05, 5.97604e-05, 5.976056e-05, 
    5.976063e-05, 5.976069e-05, 5.976084e-05, 5.976074e-05, 5.976078e-05, 
    5.976068e-05, 5.976062e-05, 5.976065e-05, 5.976046e-05, 5.976054e-05, 
    5.976015e-05, 5.976032e-05, 5.975989e-05, 5.975999e-05, 5.975987e-05, 
    5.975993e-05, 5.975982e-05, 5.975992e-05, 5.975975e-05, 5.975971e-05, 
    5.975974e-05, 5.975964e-05, 5.975992e-05, 5.975981e-05, 5.976065e-05, 
    5.976065e-05, 5.976062e-05, 5.976072e-05, 5.976073e-05, 5.976082e-05, 
    5.976074e-05, 5.976071e-05, 5.976062e-05, 5.976056e-05, 5.976051e-05, 
    5.97604e-05, 5.976028e-05, 5.976011e-05, 5.975999e-05, 5.97599e-05, 
    5.975995e-05, 5.975991e-05, 5.975996e-05, 5.975998e-05, 5.975972e-05, 
    5.975987e-05, 5.975965e-05, 5.975966e-05, 5.975976e-05, 5.975966e-05, 
    5.976064e-05, 5.976067e-05, 5.976077e-05, 5.976069e-05, 5.976083e-05, 
    5.976075e-05, 5.976071e-05, 5.976054e-05, 5.97605e-05, 5.976046e-05, 
    5.976039e-05, 5.97603e-05, 5.976014e-05, 5.976e-05, 5.975988e-05, 
    5.975989e-05, 5.975988e-05, 5.975986e-05, 5.975993e-05, 5.975985e-05, 
    5.975983e-05, 5.975987e-05, 5.975966e-05, 5.975972e-05, 5.975966e-05, 
    5.97597e-05, 5.976066e-05, 5.976062e-05, 5.976064e-05, 5.976059e-05, 
    5.976063e-05, 5.976047e-05, 5.976043e-05, 5.976022e-05, 5.97603e-05, 
    5.976016e-05, 5.976029e-05, 5.976027e-05, 5.976016e-05, 5.976028e-05, 
    5.976001e-05, 5.976019e-05, 5.975986e-05, 5.976004e-05, 5.975984e-05, 
    5.975988e-05, 5.975982e-05, 5.975977e-05, 5.975971e-05, 5.975959e-05, 
    5.975961e-05, 5.975951e-05, 5.976054e-05, 5.976048e-05, 5.976049e-05, 
    5.976042e-05, 5.976037e-05, 5.976027e-05, 5.97601e-05, 5.976016e-05, 
    5.976005e-05, 5.976003e-05, 5.97602e-05, 5.97601e-05, 5.976044e-05, 
    5.976038e-05, 5.976042e-05, 5.976054e-05, 5.976015e-05, 5.976035e-05, 
    5.975998e-05, 5.976009e-05, 5.975978e-05, 5.975994e-05, 5.975963e-05, 
    5.97595e-05, 5.975938e-05, 5.975923e-05, 5.976045e-05, 5.976049e-05, 
    5.976042e-05, 5.976031e-05, 5.976021e-05, 5.976008e-05, 5.976007e-05, 
    5.976005e-05, 5.975999e-05, 5.975993e-05, 5.976004e-05, 5.975992e-05, 
    5.976037e-05, 5.976014e-05, 5.976051e-05, 5.976039e-05, 5.976032e-05, 
    5.976035e-05, 5.976017e-05, 5.976013e-05, 5.975996e-05, 5.976005e-05, 
    5.975953e-05, 5.975976e-05, 5.975912e-05, 5.97593e-05, 5.97605e-05, 
    5.976045e-05, 5.976025e-05, 5.976034e-05, 5.976008e-05, 5.976001e-05, 
    5.975996e-05, 5.975989e-05, 5.975988e-05, 5.975984e-05, 5.975991e-05, 
    5.975984e-05, 5.976008e-05, 5.975998e-05, 5.976027e-05, 5.97602e-05, 
    5.976023e-05, 5.976027e-05, 5.976016e-05, 5.976004e-05, 5.976003e-05, 
    5.976e-05, 5.975989e-05, 5.976007e-05, 5.97595e-05, 5.975986e-05, 
    5.976039e-05, 5.976028e-05, 5.976026e-05, 5.97603e-05, 5.976002e-05, 
    5.976012e-05, 5.975984e-05, 5.975992e-05, 5.975979e-05, 5.975986e-05, 
    5.975986e-05, 5.975994e-05, 5.975999e-05, 5.976012e-05, 5.976022e-05, 
    5.97603e-05, 5.976028e-05, 5.976019e-05, 5.976003e-05, 5.975988e-05, 
    5.975991e-05, 5.97598e-05, 5.97601e-05, 5.975997e-05, 5.976002e-05, 
    5.97599e-05, 5.976017e-05, 5.975994e-05, 5.976023e-05, 5.97602e-05, 
    5.976012e-05, 5.975996e-05, 5.975993e-05, 5.975989e-05, 5.975991e-05, 
    5.976003e-05, 5.976004e-05, 5.976012e-05, 5.976015e-05, 5.976021e-05, 
    5.976026e-05, 5.976021e-05, 5.976016e-05, 5.976003e-05, 5.97599e-05, 
    5.975977e-05, 5.975974e-05, 5.975958e-05, 5.975971e-05, 5.97595e-05, 
    5.975968e-05, 5.975937e-05, 5.975992e-05, 5.975968e-05, 5.976012e-05, 
    5.976007e-05, 5.975999e-05, 5.975979e-05, 5.97599e-05, 5.975978e-05, 
    5.976004e-05, 5.976019e-05, 5.976022e-05, 5.976029e-05, 5.976022e-05, 
    5.976023e-05, 5.976016e-05, 5.976018e-05, 5.976002e-05, 5.976011e-05, 
    5.975986e-05, 5.975978e-05, 5.975952e-05, 5.975937e-05, 5.975921e-05, 
    5.975914e-05, 5.975912e-05, 5.975911e-05 ;

 TOTLITN =
  1.375895e-06, 1.375891e-06, 1.375892e-06, 1.375888e-06, 1.37589e-06, 
    1.375888e-06, 1.375894e-06, 1.375891e-06, 1.375893e-06, 1.375894e-06, 
    1.375882e-06, 1.375888e-06, 1.375876e-06, 1.375879e-06, 1.37587e-06, 
    1.375876e-06, 1.375868e-06, 1.37587e-06, 1.375865e-06, 1.375867e-06, 
    1.375861e-06, 1.375865e-06, 1.375858e-06, 1.375862e-06, 1.375861e-06, 
    1.375865e-06, 1.375887e-06, 1.375883e-06, 1.375887e-06, 1.375887e-06, 
    1.375887e-06, 1.37589e-06, 1.375892e-06, 1.375895e-06, 1.375894e-06, 
    1.375892e-06, 1.375886e-06, 1.375888e-06, 1.375883e-06, 1.375883e-06, 
    1.375878e-06, 1.37588e-06, 1.375871e-06, 1.375874e-06, 1.375867e-06, 
    1.375868e-06, 1.375867e-06, 1.375867e-06, 1.375867e-06, 1.375869e-06, 
    1.375868e-06, 1.375871e-06, 1.37588e-06, 1.375877e-06, 1.375886e-06, 
    1.375891e-06, 1.375894e-06, 1.375896e-06, 1.375896e-06, 1.375895e-06, 
    1.375892e-06, 1.375889e-06, 1.375887e-06, 1.375885e-06, 1.375883e-06, 
    1.375879e-06, 1.375876e-06, 1.375871e-06, 1.375872e-06, 1.37587e-06, 
    1.375869e-06, 1.375866e-06, 1.375866e-06, 1.375865e-06, 1.37587e-06, 
    1.375867e-06, 1.375872e-06, 1.375871e-06, 1.375883e-06, 1.375888e-06, 
    1.37589e-06, 1.375891e-06, 1.375896e-06, 1.375893e-06, 1.375894e-06, 
    1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375885e-06, 1.375887e-06, 
    1.375876e-06, 1.375881e-06, 1.375869e-06, 1.375872e-06, 1.375868e-06, 
    1.37587e-06, 1.375867e-06, 1.37587e-06, 1.375865e-06, 1.375864e-06, 
    1.375864e-06, 1.375862e-06, 1.37587e-06, 1.375867e-06, 1.37589e-06, 
    1.37589e-06, 1.375889e-06, 1.375892e-06, 1.375892e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375889e-06, 1.375888e-06, 1.375886e-06, 
    1.375883e-06, 1.37588e-06, 1.375875e-06, 1.375871e-06, 1.375869e-06, 
    1.375871e-06, 1.375869e-06, 1.375871e-06, 1.375871e-06, 1.375864e-06, 
    1.375868e-06, 1.375862e-06, 1.375862e-06, 1.375865e-06, 1.375862e-06, 
    1.37589e-06, 1.375891e-06, 1.375894e-06, 1.375891e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375887e-06, 1.375886e-06, 1.375885e-06, 
    1.375883e-06, 1.37588e-06, 1.375876e-06, 1.375872e-06, 1.375868e-06, 
    1.375869e-06, 1.375869e-06, 1.375868e-06, 1.37587e-06, 1.375868e-06, 
    1.375867e-06, 1.375868e-06, 1.375862e-06, 1.375864e-06, 1.375862e-06, 
    1.375863e-06, 1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375889e-06, 
    1.375889e-06, 1.375885e-06, 1.375884e-06, 1.375878e-06, 1.37588e-06, 
    1.375876e-06, 1.37588e-06, 1.375879e-06, 1.375876e-06, 1.37588e-06, 
    1.375872e-06, 1.375877e-06, 1.375868e-06, 1.375873e-06, 1.375868e-06, 
    1.375868e-06, 1.375867e-06, 1.375865e-06, 1.375864e-06, 1.37586e-06, 
    1.375861e-06, 1.375858e-06, 1.375887e-06, 1.375885e-06, 1.375886e-06, 
    1.375884e-06, 1.375882e-06, 1.375879e-06, 1.375875e-06, 1.375877e-06, 
    1.375873e-06, 1.375873e-06, 1.375878e-06, 1.375875e-06, 1.375884e-06, 
    1.375883e-06, 1.375884e-06, 1.375887e-06, 1.375876e-06, 1.375882e-06, 
    1.375871e-06, 1.375874e-06, 1.375866e-06, 1.37587e-06, 1.375861e-06, 
    1.375858e-06, 1.375854e-06, 1.37585e-06, 1.375884e-06, 1.375886e-06, 
    1.375883e-06, 1.375881e-06, 1.375878e-06, 1.375874e-06, 1.375874e-06, 
    1.375873e-06, 1.375871e-06, 1.37587e-06, 1.375873e-06, 1.37587e-06, 
    1.375882e-06, 1.375876e-06, 1.375886e-06, 1.375883e-06, 1.375881e-06, 
    1.375882e-06, 1.375877e-06, 1.375876e-06, 1.375871e-06, 1.375873e-06, 
    1.375859e-06, 1.375865e-06, 1.375847e-06, 1.375852e-06, 1.375886e-06, 
    1.375884e-06, 1.375879e-06, 1.375882e-06, 1.375874e-06, 1.375872e-06, 
    1.375871e-06, 1.375869e-06, 1.375868e-06, 1.375867e-06, 1.375869e-06, 
    1.375867e-06, 1.375874e-06, 1.375871e-06, 1.375879e-06, 1.375878e-06, 
    1.375878e-06, 1.375879e-06, 1.375876e-06, 1.375873e-06, 1.375873e-06, 
    1.375872e-06, 1.375869e-06, 1.375874e-06, 1.375858e-06, 1.375868e-06, 
    1.375883e-06, 1.37588e-06, 1.375879e-06, 1.37588e-06, 1.375872e-06, 
    1.375875e-06, 1.375867e-06, 1.375869e-06, 1.375866e-06, 1.375868e-06, 
    1.375868e-06, 1.37587e-06, 1.375872e-06, 1.375875e-06, 1.375878e-06, 
    1.37588e-06, 1.37588e-06, 1.375877e-06, 1.375873e-06, 1.375868e-06, 
    1.375869e-06, 1.375866e-06, 1.375875e-06, 1.375871e-06, 1.375872e-06, 
    1.375869e-06, 1.375877e-06, 1.37587e-06, 1.375878e-06, 1.375878e-06, 
    1.375875e-06, 1.375871e-06, 1.37587e-06, 1.375869e-06, 1.375869e-06, 
    1.375873e-06, 1.375873e-06, 1.375875e-06, 1.375876e-06, 1.375878e-06, 
    1.375879e-06, 1.375878e-06, 1.375876e-06, 1.375873e-06, 1.375869e-06, 
    1.375865e-06, 1.375864e-06, 1.37586e-06, 1.375864e-06, 1.375858e-06, 
    1.375863e-06, 1.375854e-06, 1.37587e-06, 1.375863e-06, 1.375875e-06, 
    1.375874e-06, 1.375872e-06, 1.375866e-06, 1.375869e-06, 1.375866e-06, 
    1.375873e-06, 1.375877e-06, 1.375878e-06, 1.37588e-06, 1.375878e-06, 
    1.375878e-06, 1.375876e-06, 1.375877e-06, 1.375872e-06, 1.375875e-06, 
    1.375868e-06, 1.375866e-06, 1.375858e-06, 1.375854e-06, 1.37585e-06, 
    1.375848e-06, 1.375847e-06, 1.375847e-06 ;

 TOTLITN_1m =
  1.375895e-06, 1.375891e-06, 1.375892e-06, 1.375888e-06, 1.37589e-06, 
    1.375888e-06, 1.375894e-06, 1.375891e-06, 1.375893e-06, 1.375894e-06, 
    1.375882e-06, 1.375888e-06, 1.375876e-06, 1.375879e-06, 1.37587e-06, 
    1.375876e-06, 1.375868e-06, 1.37587e-06, 1.375865e-06, 1.375867e-06, 
    1.375861e-06, 1.375865e-06, 1.375858e-06, 1.375862e-06, 1.375861e-06, 
    1.375865e-06, 1.375887e-06, 1.375883e-06, 1.375887e-06, 1.375887e-06, 
    1.375887e-06, 1.37589e-06, 1.375892e-06, 1.375895e-06, 1.375894e-06, 
    1.375892e-06, 1.375886e-06, 1.375888e-06, 1.375883e-06, 1.375883e-06, 
    1.375878e-06, 1.37588e-06, 1.375871e-06, 1.375874e-06, 1.375867e-06, 
    1.375868e-06, 1.375867e-06, 1.375867e-06, 1.375867e-06, 1.375869e-06, 
    1.375868e-06, 1.375871e-06, 1.37588e-06, 1.375877e-06, 1.375886e-06, 
    1.375891e-06, 1.375894e-06, 1.375896e-06, 1.375896e-06, 1.375895e-06, 
    1.375892e-06, 1.375889e-06, 1.375887e-06, 1.375885e-06, 1.375883e-06, 
    1.375879e-06, 1.375876e-06, 1.375871e-06, 1.375872e-06, 1.37587e-06, 
    1.375869e-06, 1.375866e-06, 1.375866e-06, 1.375865e-06, 1.37587e-06, 
    1.375867e-06, 1.375872e-06, 1.375871e-06, 1.375883e-06, 1.375888e-06, 
    1.37589e-06, 1.375891e-06, 1.375896e-06, 1.375893e-06, 1.375894e-06, 
    1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375885e-06, 1.375887e-06, 
    1.375876e-06, 1.375881e-06, 1.375869e-06, 1.375872e-06, 1.375868e-06, 
    1.37587e-06, 1.375867e-06, 1.37587e-06, 1.375865e-06, 1.375864e-06, 
    1.375864e-06, 1.375862e-06, 1.37587e-06, 1.375867e-06, 1.37589e-06, 
    1.37589e-06, 1.375889e-06, 1.375892e-06, 1.375892e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375889e-06, 1.375888e-06, 1.375886e-06, 
    1.375883e-06, 1.37588e-06, 1.375875e-06, 1.375871e-06, 1.375869e-06, 
    1.375871e-06, 1.375869e-06, 1.375871e-06, 1.375871e-06, 1.375864e-06, 
    1.375868e-06, 1.375862e-06, 1.375862e-06, 1.375865e-06, 1.375862e-06, 
    1.37589e-06, 1.375891e-06, 1.375894e-06, 1.375891e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375887e-06, 1.375886e-06, 1.375885e-06, 
    1.375883e-06, 1.37588e-06, 1.375876e-06, 1.375872e-06, 1.375868e-06, 
    1.375869e-06, 1.375869e-06, 1.375868e-06, 1.37587e-06, 1.375868e-06, 
    1.375867e-06, 1.375868e-06, 1.375862e-06, 1.375864e-06, 1.375862e-06, 
    1.375863e-06, 1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375889e-06, 
    1.375889e-06, 1.375885e-06, 1.375884e-06, 1.375878e-06, 1.37588e-06, 
    1.375876e-06, 1.37588e-06, 1.375879e-06, 1.375876e-06, 1.37588e-06, 
    1.375872e-06, 1.375877e-06, 1.375868e-06, 1.375873e-06, 1.375868e-06, 
    1.375868e-06, 1.375867e-06, 1.375865e-06, 1.375864e-06, 1.37586e-06, 
    1.375861e-06, 1.375858e-06, 1.375887e-06, 1.375885e-06, 1.375886e-06, 
    1.375884e-06, 1.375882e-06, 1.375879e-06, 1.375875e-06, 1.375877e-06, 
    1.375873e-06, 1.375873e-06, 1.375878e-06, 1.375875e-06, 1.375884e-06, 
    1.375883e-06, 1.375884e-06, 1.375887e-06, 1.375876e-06, 1.375882e-06, 
    1.375871e-06, 1.375874e-06, 1.375866e-06, 1.37587e-06, 1.375861e-06, 
    1.375858e-06, 1.375854e-06, 1.37585e-06, 1.375884e-06, 1.375886e-06, 
    1.375883e-06, 1.375881e-06, 1.375878e-06, 1.375874e-06, 1.375874e-06, 
    1.375873e-06, 1.375871e-06, 1.37587e-06, 1.375873e-06, 1.37587e-06, 
    1.375882e-06, 1.375876e-06, 1.375886e-06, 1.375883e-06, 1.375881e-06, 
    1.375882e-06, 1.375877e-06, 1.375876e-06, 1.375871e-06, 1.375873e-06, 
    1.375859e-06, 1.375865e-06, 1.375847e-06, 1.375852e-06, 1.375886e-06, 
    1.375884e-06, 1.375879e-06, 1.375882e-06, 1.375874e-06, 1.375872e-06, 
    1.375871e-06, 1.375869e-06, 1.375868e-06, 1.375867e-06, 1.375869e-06, 
    1.375867e-06, 1.375874e-06, 1.375871e-06, 1.375879e-06, 1.375878e-06, 
    1.375878e-06, 1.375879e-06, 1.375876e-06, 1.375873e-06, 1.375873e-06, 
    1.375872e-06, 1.375869e-06, 1.375874e-06, 1.375858e-06, 1.375868e-06, 
    1.375883e-06, 1.37588e-06, 1.375879e-06, 1.37588e-06, 1.375872e-06, 
    1.375875e-06, 1.375867e-06, 1.375869e-06, 1.375866e-06, 1.375868e-06, 
    1.375868e-06, 1.37587e-06, 1.375872e-06, 1.375875e-06, 1.375878e-06, 
    1.37588e-06, 1.37588e-06, 1.375877e-06, 1.375873e-06, 1.375868e-06, 
    1.375869e-06, 1.375866e-06, 1.375875e-06, 1.375871e-06, 1.375872e-06, 
    1.375869e-06, 1.375877e-06, 1.37587e-06, 1.375878e-06, 1.375878e-06, 
    1.375875e-06, 1.375871e-06, 1.37587e-06, 1.375869e-06, 1.375869e-06, 
    1.375873e-06, 1.375873e-06, 1.375875e-06, 1.375876e-06, 1.375878e-06, 
    1.375879e-06, 1.375878e-06, 1.375876e-06, 1.375873e-06, 1.375869e-06, 
    1.375865e-06, 1.375864e-06, 1.37586e-06, 1.375864e-06, 1.375858e-06, 
    1.375863e-06, 1.375854e-06, 1.37587e-06, 1.375863e-06, 1.375875e-06, 
    1.375874e-06, 1.375872e-06, 1.375866e-06, 1.375869e-06, 1.375866e-06, 
    1.375873e-06, 1.375877e-06, 1.375878e-06, 1.37588e-06, 1.375878e-06, 
    1.375878e-06, 1.375876e-06, 1.375877e-06, 1.375872e-06, 1.375875e-06, 
    1.375868e-06, 1.375866e-06, 1.375858e-06, 1.375854e-06, 1.37585e-06, 
    1.375848e-06, 1.375847e-06, 1.375847e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34412, 17.34411, 17.34411, 17.3441, 17.34411, 17.3441, 17.34412, 
    17.34411, 17.34411, 17.34412, 17.34409, 17.3441, 17.34407, 17.34408, 
    17.34406, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34404, 
    17.34405, 17.34403, 17.34404, 17.34404, 17.34405, 17.3441, 17.34409, 
    17.3441, 17.3441, 17.3441, 17.34411, 17.34411, 17.34412, 17.34412, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34409, 
    17.34406, 17.34407, 17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 
    17.34406, 17.34406, 17.34406, 17.34408, 17.34408, 17.3441, 17.34411, 
    17.34412, 17.34412, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 
    17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34406, 17.34409, 17.3441, 17.34411, 17.34411, 17.34412, 17.34411, 
    17.34412, 17.34411, 17.34411, 17.34411, 17.3441, 17.3441, 17.34407, 
    17.34409, 17.34406, 17.34406, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34404, 17.34405, 17.34404, 17.34406, 17.34405, 17.34411, 
    17.34411, 17.34411, 17.34411, 17.34411, 17.34412, 17.34411, 17.34411, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34406, 17.34406, 17.34406, 17.34406, 17.34404, 17.34406, 
    17.34404, 17.34404, 17.34405, 17.34404, 17.34411, 17.34411, 17.34412, 
    17.34411, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 17.3441, 
    17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34406, 17.34404, 17.34404, 
    17.34404, 17.34404, 17.34411, 17.34411, 17.34411, 17.3441, 17.34411, 
    17.3441, 17.34409, 17.34408, 17.34408, 17.34407, 17.34408, 17.34408, 
    17.34407, 17.34408, 17.34406, 17.34408, 17.34405, 17.34407, 17.34405, 
    17.34406, 17.34405, 17.34405, 17.34404, 17.34403, 17.34404, 17.34403, 
    17.3441, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34407, 
    17.34407, 17.34407, 17.34406, 17.34408, 17.34407, 17.34409, 17.34409, 
    17.34409, 17.3441, 17.34407, 17.34409, 17.34406, 17.34407, 17.34405, 
    17.34406, 17.34404, 17.34403, 17.34402, 17.34401, 17.3441, 17.3441, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34407, 17.34407, 17.34406, 
    17.34406, 17.34407, 17.34406, 17.34409, 17.34407, 17.3441, 17.34409, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.344, 17.34402, 17.3441, 17.3441, 17.34408, 17.34409, 
    17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34407, 17.34406, 17.34408, 17.34408, 17.34408, 17.34408, 
    17.34407, 17.34407, 17.34407, 17.34406, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.34409, 17.34408, 17.34408, 17.34408, 17.34406, 17.34407, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34406, 
    17.34407, 17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34405, 17.34407, 17.34406, 17.34406, 17.34406, 17.34408, 
    17.34406, 17.34408, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34406, 17.34407, 17.34407, 17.34407, 17.34408, 17.34408, 
    17.34408, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34403, 
    17.34404, 17.34403, 17.34404, 17.34402, 17.34406, 17.34404, 17.34407, 
    17.34407, 17.34406, 17.34405, 17.34406, 17.34405, 17.34407, 17.34408, 
    17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34408, 17.34406, 
    17.34407, 17.34405, 17.34405, 17.34403, 17.34402, 17.34401, 17.344, 
    17.344, 17.344 ;

 TOTSOMC_1m =
  17.34412, 17.34411, 17.34411, 17.3441, 17.34411, 17.3441, 17.34412, 
    17.34411, 17.34411, 17.34412, 17.34409, 17.3441, 17.34407, 17.34408, 
    17.34406, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34404, 
    17.34405, 17.34403, 17.34404, 17.34404, 17.34405, 17.3441, 17.34409, 
    17.3441, 17.3441, 17.3441, 17.34411, 17.34411, 17.34412, 17.34412, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34409, 
    17.34406, 17.34407, 17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 
    17.34406, 17.34406, 17.34406, 17.34408, 17.34408, 17.3441, 17.34411, 
    17.34412, 17.34412, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 
    17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34406, 17.34409, 17.3441, 17.34411, 17.34411, 17.34412, 17.34411, 
    17.34412, 17.34411, 17.34411, 17.34411, 17.3441, 17.3441, 17.34407, 
    17.34409, 17.34406, 17.34406, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34404, 17.34405, 17.34404, 17.34406, 17.34405, 17.34411, 
    17.34411, 17.34411, 17.34411, 17.34411, 17.34412, 17.34411, 17.34411, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34406, 17.34406, 17.34406, 17.34406, 17.34404, 17.34406, 
    17.34404, 17.34404, 17.34405, 17.34404, 17.34411, 17.34411, 17.34412, 
    17.34411, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 17.3441, 
    17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34406, 17.34404, 17.34404, 
    17.34404, 17.34404, 17.34411, 17.34411, 17.34411, 17.3441, 17.34411, 
    17.3441, 17.34409, 17.34408, 17.34408, 17.34407, 17.34408, 17.34408, 
    17.34407, 17.34408, 17.34406, 17.34408, 17.34405, 17.34407, 17.34405, 
    17.34406, 17.34405, 17.34405, 17.34404, 17.34403, 17.34404, 17.34403, 
    17.3441, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34407, 
    17.34407, 17.34407, 17.34406, 17.34408, 17.34407, 17.34409, 17.34409, 
    17.34409, 17.3441, 17.34407, 17.34409, 17.34406, 17.34407, 17.34405, 
    17.34406, 17.34404, 17.34403, 17.34402, 17.34401, 17.3441, 17.3441, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34407, 17.34407, 17.34406, 
    17.34406, 17.34407, 17.34406, 17.34409, 17.34407, 17.3441, 17.34409, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.344, 17.34402, 17.3441, 17.3441, 17.34408, 17.34409, 
    17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34407, 17.34406, 17.34408, 17.34408, 17.34408, 17.34408, 
    17.34407, 17.34407, 17.34407, 17.34406, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.34409, 17.34408, 17.34408, 17.34408, 17.34406, 17.34407, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34406, 
    17.34407, 17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34405, 17.34407, 17.34406, 17.34406, 17.34406, 17.34408, 
    17.34406, 17.34408, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34406, 17.34407, 17.34407, 17.34407, 17.34408, 17.34408, 
    17.34408, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34403, 
    17.34404, 17.34403, 17.34404, 17.34402, 17.34406, 17.34404, 17.34407, 
    17.34407, 17.34406, 17.34405, 17.34406, 17.34405, 17.34407, 17.34408, 
    17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34408, 17.34406, 
    17.34407, 17.34405, 17.34405, 17.34403, 17.34402, 17.34401, 17.344, 
    17.344, 17.344 ;

 TOTSOMN =
  1.773689, 1.773688, 1.773688, 1.773687, 1.773688, 1.773687, 1.773689, 
    1.773688, 1.773689, 1.773689, 1.773685, 1.773687, 1.773683, 1.773684, 
    1.773681, 1.773683, 1.77368, 1.773681, 1.773679, 1.773679, 1.773677, 
    1.773679, 1.773676, 1.773678, 1.773678, 1.773679, 1.773687, 1.773685, 
    1.773687, 1.773686, 1.773687, 1.773688, 1.773688, 1.773689, 1.773689, 
    1.773688, 1.773686, 1.773687, 1.773685, 1.773685, 1.773683, 1.773684, 
    1.773681, 1.773682, 1.773679, 1.77368, 1.773679, 1.77368, 1.773679, 
    1.77368, 1.77368, 1.773681, 1.773684, 1.773683, 1.773686, 1.773688, 
    1.773689, 1.77369, 1.77369, 1.77369, 1.773688, 1.773687, 1.773686, 
    1.773686, 1.773685, 1.773684, 1.773683, 1.773681, 1.773681, 1.773681, 
    1.77368, 1.773679, 1.773679, 1.773679, 1.773681, 1.77368, 1.773682, 
    1.773681, 1.773685, 1.773687, 1.773687, 1.773688, 1.77369, 1.773689, 
    1.773689, 1.773688, 1.773687, 1.773688, 1.773686, 1.773687, 1.773683, 
    1.773685, 1.77368, 1.773681, 1.77368, 1.773681, 1.773679, 1.773681, 
    1.773679, 1.773678, 1.773679, 1.773678, 1.773681, 1.773679, 1.773688, 
    1.773688, 1.773687, 1.773688, 1.773689, 1.773689, 1.773689, 1.773688, 
    1.773687, 1.773687, 1.773686, 1.773685, 1.773684, 1.773682, 1.773681, 
    1.77368, 1.773681, 1.77368, 1.773681, 1.773681, 1.773679, 1.77368, 
    1.773678, 1.773678, 1.773679, 1.773678, 1.773688, 1.773688, 1.773689, 
    1.773688, 1.77369, 1.773689, 1.773688, 1.773687, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773681, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773681, 1.77368, 1.77368, 1.77368, 1.773678, 1.773679, 
    1.773678, 1.773678, 1.773688, 1.773687, 1.773688, 1.773687, 1.773687, 
    1.773686, 1.773686, 1.773683, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773684, 1.773681, 1.773683, 1.77368, 1.773682, 1.77368, 
    1.77368, 1.77368, 1.773679, 1.773678, 1.773677, 1.773677, 1.773677, 
    1.773687, 1.773686, 1.773686, 1.773685, 1.773685, 1.773684, 1.773682, 
    1.773683, 1.773682, 1.773682, 1.773683, 1.773682, 1.773686, 1.773685, 
    1.773685, 1.773687, 1.773683, 1.773685, 1.773681, 1.773682, 1.773679, 
    1.773681, 1.773678, 1.773676, 1.773675, 1.773674, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773682, 1.773682, 1.773682, 1.773681, 
    1.773681, 1.773682, 1.773681, 1.773685, 1.773683, 1.773686, 1.773685, 
    1.773684, 1.773685, 1.773683, 1.773683, 1.773681, 1.773682, 1.773677, 
    1.773679, 1.773673, 1.773674, 1.773686, 1.773686, 1.773684, 1.773685, 
    1.773682, 1.773681, 1.773681, 1.77368, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773682, 1.773681, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773682, 1.773682, 1.773681, 1.77368, 1.773682, 1.773676, 
    1.77368, 1.773685, 1.773684, 1.773684, 1.773684, 1.773682, 1.773682, 
    1.77368, 1.773681, 1.773679, 1.77368, 1.77368, 1.773681, 1.773681, 
    1.773682, 1.773683, 1.773684, 1.773684, 1.773683, 1.773682, 1.77368, 
    1.77368, 1.773679, 1.773682, 1.773681, 1.773682, 1.77368, 1.773683, 
    1.773681, 1.773684, 1.773683, 1.773683, 1.773681, 1.773681, 1.77368, 
    1.77368, 1.773682, 1.773682, 1.773683, 1.773683, 1.773683, 1.773684, 
    1.773683, 1.773683, 1.773682, 1.77368, 1.773679, 1.773679, 1.773677, 
    1.773678, 1.773676, 1.773678, 1.773675, 1.773681, 1.773678, 1.773682, 
    1.773682, 1.773681, 1.773679, 1.77368, 1.773679, 1.773682, 1.773683, 
    1.773684, 1.773684, 1.773684, 1.773684, 1.773683, 1.773683, 1.773682, 
    1.773682, 1.77368, 1.773679, 1.773677, 1.773675, 1.773674, 1.773673, 
    1.773673, 1.773673 ;

 TOTSOMN_1m =
  1.773689, 1.773688, 1.773688, 1.773687, 1.773688, 1.773687, 1.773689, 
    1.773688, 1.773689, 1.773689, 1.773685, 1.773687, 1.773683, 1.773684, 
    1.773681, 1.773683, 1.77368, 1.773681, 1.773679, 1.773679, 1.773677, 
    1.773679, 1.773676, 1.773678, 1.773678, 1.773679, 1.773687, 1.773685, 
    1.773687, 1.773686, 1.773687, 1.773688, 1.773688, 1.773689, 1.773689, 
    1.773688, 1.773686, 1.773687, 1.773685, 1.773685, 1.773683, 1.773684, 
    1.773681, 1.773682, 1.773679, 1.77368, 1.773679, 1.77368, 1.773679, 
    1.77368, 1.77368, 1.773681, 1.773684, 1.773683, 1.773686, 1.773688, 
    1.773689, 1.77369, 1.77369, 1.77369, 1.773688, 1.773687, 1.773686, 
    1.773686, 1.773685, 1.773684, 1.773683, 1.773681, 1.773681, 1.773681, 
    1.77368, 1.773679, 1.773679, 1.773679, 1.773681, 1.77368, 1.773682, 
    1.773681, 1.773685, 1.773687, 1.773687, 1.773688, 1.77369, 1.773689, 
    1.773689, 1.773688, 1.773687, 1.773688, 1.773686, 1.773687, 1.773683, 
    1.773685, 1.77368, 1.773681, 1.77368, 1.773681, 1.773679, 1.773681, 
    1.773679, 1.773678, 1.773679, 1.773678, 1.773681, 1.773679, 1.773688, 
    1.773688, 1.773687, 1.773688, 1.773689, 1.773689, 1.773689, 1.773688, 
    1.773687, 1.773687, 1.773686, 1.773685, 1.773684, 1.773682, 1.773681, 
    1.77368, 1.773681, 1.77368, 1.773681, 1.773681, 1.773679, 1.77368, 
    1.773678, 1.773678, 1.773679, 1.773678, 1.773688, 1.773688, 1.773689, 
    1.773688, 1.77369, 1.773689, 1.773688, 1.773687, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773681, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773681, 1.77368, 1.77368, 1.77368, 1.773678, 1.773679, 
    1.773678, 1.773678, 1.773688, 1.773687, 1.773688, 1.773687, 1.773687, 
    1.773686, 1.773686, 1.773683, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773684, 1.773681, 1.773683, 1.77368, 1.773682, 1.77368, 
    1.77368, 1.77368, 1.773679, 1.773678, 1.773677, 1.773677, 1.773677, 
    1.773687, 1.773686, 1.773686, 1.773685, 1.773685, 1.773684, 1.773682, 
    1.773683, 1.773682, 1.773682, 1.773683, 1.773682, 1.773686, 1.773685, 
    1.773685, 1.773687, 1.773683, 1.773685, 1.773681, 1.773682, 1.773679, 
    1.773681, 1.773678, 1.773676, 1.773675, 1.773674, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773682, 1.773682, 1.773682, 1.773681, 
    1.773681, 1.773682, 1.773681, 1.773685, 1.773683, 1.773686, 1.773685, 
    1.773684, 1.773685, 1.773683, 1.773683, 1.773681, 1.773682, 1.773677, 
    1.773679, 1.773673, 1.773674, 1.773686, 1.773686, 1.773684, 1.773685, 
    1.773682, 1.773681, 1.773681, 1.77368, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773682, 1.773681, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773682, 1.773682, 1.773681, 1.77368, 1.773682, 1.773676, 
    1.77368, 1.773685, 1.773684, 1.773684, 1.773684, 1.773682, 1.773682, 
    1.77368, 1.773681, 1.773679, 1.77368, 1.77368, 1.773681, 1.773681, 
    1.773682, 1.773683, 1.773684, 1.773684, 1.773683, 1.773682, 1.77368, 
    1.77368, 1.773679, 1.773682, 1.773681, 1.773682, 1.77368, 1.773683, 
    1.773681, 1.773684, 1.773683, 1.773683, 1.773681, 1.773681, 1.77368, 
    1.77368, 1.773682, 1.773682, 1.773683, 1.773683, 1.773683, 1.773684, 
    1.773683, 1.773683, 1.773682, 1.77368, 1.773679, 1.773679, 1.773677, 
    1.773678, 1.773676, 1.773678, 1.773675, 1.773681, 1.773678, 1.773682, 
    1.773682, 1.773681, 1.773679, 1.77368, 1.773679, 1.773682, 1.773683, 
    1.773684, 1.773684, 1.773684, 1.773684, 1.773683, 1.773683, 1.773682, 
    1.773682, 1.77368, 1.773679, 1.773677, 1.773675, 1.773674, 1.773673, 
    1.773673, 1.773673 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.992, 249.9922, 249.9922, 249.9924, 249.9922, 249.9924, 249.992, 
    249.9922, 249.9921, 249.992, 249.9927, 249.9924, 249.9931, 249.9929, 
    249.9935, 249.9931, 249.9935, 249.9935, 249.9937, 249.9937, 249.994, 
    249.9938, 249.9942, 249.9939, 249.994, 249.9938, 249.9924, 249.9927, 
    249.9924, 249.9925, 249.9924, 249.9922, 249.9922, 249.992, 249.992, 
    249.9921, 249.9925, 249.9924, 249.9927, 249.9926, 249.993, 249.9928, 
    249.9934, 249.9932, 249.9937, 249.9935, 249.9937, 249.9936, 249.9937, 
    249.9935, 249.9936, 249.9934, 249.9929, 249.993, 249.9925, 249.9922, 
    249.992, 249.9919, 249.9919, 249.9919, 249.9921, 249.9923, 249.9925, 
    249.9926, 249.9926, 249.9929, 249.9931, 249.9934, 249.9933, 249.9934, 
    249.9935, 249.9937, 249.9937, 249.9937, 249.9934, 249.9936, 249.9933, 
    249.9934, 249.9927, 249.9924, 249.9923, 249.9922, 249.9919, 249.9921, 
    249.992, 249.9922, 249.9923, 249.9922, 249.9926, 249.9924, 249.9931, 
    249.9928, 249.9935, 249.9933, 249.9936, 249.9935, 249.9937, 249.9935, 
    249.9938, 249.9938, 249.9938, 249.994, 249.9935, 249.9937, 249.9922, 
    249.9922, 249.9923, 249.9921, 249.9921, 249.992, 249.9921, 249.9922, 
    249.9923, 249.9924, 249.9925, 249.9927, 249.9929, 249.9931, 249.9934, 
    249.9935, 249.9934, 249.9935, 249.9934, 249.9934, 249.9938, 249.9936, 
    249.9939, 249.9939, 249.9937, 249.9939, 249.9923, 249.9922, 249.9921, 
    249.9922, 249.9919, 249.9921, 249.9921, 249.9924, 249.9925, 249.9926, 
    249.9927, 249.9928, 249.9931, 249.9933, 249.9935, 249.9935, 249.9935, 
    249.9936, 249.9935, 249.9936, 249.9936, 249.9936, 249.9939, 249.9938, 
    249.9939, 249.9939, 249.9922, 249.9923, 249.9923, 249.9923, 249.9923, 
    249.9925, 249.9926, 249.993, 249.9928, 249.9931, 249.9929, 249.9929, 
    249.9931, 249.9929, 249.9933, 249.993, 249.9936, 249.9933, 249.9936, 
    249.9935, 249.9936, 249.9937, 249.9938, 249.994, 249.994, 249.9942, 
    249.9924, 249.9925, 249.9925, 249.9926, 249.9927, 249.9929, 249.9932, 
    249.9931, 249.9933, 249.9933, 249.993, 249.9932, 249.9926, 249.9927, 
    249.9926, 249.9924, 249.9931, 249.9928, 249.9934, 249.9932, 249.9937, 
    249.9935, 249.994, 249.9942, 249.9944, 249.9946, 249.9926, 249.9925, 
    249.9926, 249.9928, 249.993, 249.9932, 249.9932, 249.9933, 249.9934, 
    249.9935, 249.9933, 249.9935, 249.9927, 249.9931, 249.9925, 249.9927, 
    249.9928, 249.9928, 249.9931, 249.9931, 249.9934, 249.9933, 249.9941, 
    249.9937, 249.9948, 249.9945, 249.9925, 249.9926, 249.9929, 249.9928, 
    249.9932, 249.9933, 249.9934, 249.9935, 249.9935, 249.9936, 249.9935, 
    249.9936, 249.9932, 249.9934, 249.9929, 249.993, 249.993, 249.9929, 
    249.9931, 249.9933, 249.9933, 249.9933, 249.9935, 249.9932, 249.9942, 
    249.9936, 249.9927, 249.9929, 249.9929, 249.9928, 249.9933, 249.9931, 
    249.9936, 249.9935, 249.9937, 249.9936, 249.9936, 249.9934, 249.9934, 
    249.9931, 249.993, 249.9928, 249.9929, 249.993, 249.9933, 249.9935, 
    249.9935, 249.9937, 249.9932, 249.9934, 249.9933, 249.9935, 249.9931, 
    249.9934, 249.993, 249.993, 249.9931, 249.9934, 249.9935, 249.9935, 
    249.9935, 249.9933, 249.9933, 249.9931, 249.9931, 249.993, 249.9929, 
    249.993, 249.9931, 249.9933, 249.9935, 249.9937, 249.9938, 249.994, 
    249.9938, 249.9942, 249.9939, 249.9944, 249.9935, 249.9939, 249.9931, 
    249.9932, 249.9934, 249.9937, 249.9935, 249.9937, 249.9933, 249.993, 
    249.993, 249.9928, 249.993, 249.993, 249.9931, 249.993, 249.9933, 
    249.9932, 249.9936, 249.9937, 249.9941, 249.9944, 249.9947, 249.9948, 
    249.9948, 249.9948 ;

 TREFMNAV_R =
  249.992, 249.9922, 249.9922, 249.9924, 249.9922, 249.9924, 249.992, 
    249.9922, 249.9921, 249.992, 249.9927, 249.9924, 249.9931, 249.9929, 
    249.9935, 249.9931, 249.9935, 249.9935, 249.9937, 249.9937, 249.994, 
    249.9938, 249.9942, 249.9939, 249.994, 249.9938, 249.9924, 249.9927, 
    249.9924, 249.9925, 249.9924, 249.9922, 249.9922, 249.992, 249.992, 
    249.9921, 249.9925, 249.9924, 249.9927, 249.9926, 249.993, 249.9928, 
    249.9934, 249.9932, 249.9937, 249.9935, 249.9937, 249.9936, 249.9937, 
    249.9935, 249.9936, 249.9934, 249.9929, 249.993, 249.9925, 249.9922, 
    249.992, 249.9919, 249.9919, 249.9919, 249.9921, 249.9923, 249.9925, 
    249.9926, 249.9926, 249.9929, 249.9931, 249.9934, 249.9933, 249.9934, 
    249.9935, 249.9937, 249.9937, 249.9937, 249.9934, 249.9936, 249.9933, 
    249.9934, 249.9927, 249.9924, 249.9923, 249.9922, 249.9919, 249.9921, 
    249.992, 249.9922, 249.9923, 249.9922, 249.9926, 249.9924, 249.9931, 
    249.9928, 249.9935, 249.9933, 249.9936, 249.9935, 249.9937, 249.9935, 
    249.9938, 249.9938, 249.9938, 249.994, 249.9935, 249.9937, 249.9922, 
    249.9922, 249.9923, 249.9921, 249.9921, 249.992, 249.9921, 249.9922, 
    249.9923, 249.9924, 249.9925, 249.9927, 249.9929, 249.9931, 249.9934, 
    249.9935, 249.9934, 249.9935, 249.9934, 249.9934, 249.9938, 249.9936, 
    249.9939, 249.9939, 249.9937, 249.9939, 249.9923, 249.9922, 249.9921, 
    249.9922, 249.9919, 249.9921, 249.9921, 249.9924, 249.9925, 249.9926, 
    249.9927, 249.9928, 249.9931, 249.9933, 249.9935, 249.9935, 249.9935, 
    249.9936, 249.9935, 249.9936, 249.9936, 249.9936, 249.9939, 249.9938, 
    249.9939, 249.9939, 249.9922, 249.9923, 249.9923, 249.9923, 249.9923, 
    249.9925, 249.9926, 249.993, 249.9928, 249.9931, 249.9929, 249.9929, 
    249.9931, 249.9929, 249.9933, 249.993, 249.9936, 249.9933, 249.9936, 
    249.9935, 249.9936, 249.9937, 249.9938, 249.994, 249.994, 249.9942, 
    249.9924, 249.9925, 249.9925, 249.9926, 249.9927, 249.9929, 249.9932, 
    249.9931, 249.9933, 249.9933, 249.993, 249.9932, 249.9926, 249.9927, 
    249.9926, 249.9924, 249.9931, 249.9928, 249.9934, 249.9932, 249.9937, 
    249.9935, 249.994, 249.9942, 249.9944, 249.9946, 249.9926, 249.9925, 
    249.9926, 249.9928, 249.993, 249.9932, 249.9932, 249.9933, 249.9934, 
    249.9935, 249.9933, 249.9935, 249.9927, 249.9931, 249.9925, 249.9927, 
    249.9928, 249.9928, 249.9931, 249.9931, 249.9934, 249.9933, 249.9941, 
    249.9937, 249.9948, 249.9945, 249.9925, 249.9926, 249.9929, 249.9928, 
    249.9932, 249.9933, 249.9934, 249.9935, 249.9935, 249.9936, 249.9935, 
    249.9936, 249.9932, 249.9934, 249.9929, 249.993, 249.993, 249.9929, 
    249.9931, 249.9933, 249.9933, 249.9933, 249.9935, 249.9932, 249.9942, 
    249.9936, 249.9927, 249.9929, 249.9929, 249.9928, 249.9933, 249.9931, 
    249.9936, 249.9935, 249.9937, 249.9936, 249.9936, 249.9934, 249.9934, 
    249.9931, 249.993, 249.9928, 249.9929, 249.993, 249.9933, 249.9935, 
    249.9935, 249.9937, 249.9932, 249.9934, 249.9933, 249.9935, 249.9931, 
    249.9934, 249.993, 249.993, 249.9931, 249.9934, 249.9935, 249.9935, 
    249.9935, 249.9933, 249.9933, 249.9931, 249.9931, 249.993, 249.9929, 
    249.993, 249.9931, 249.9933, 249.9935, 249.9937, 249.9938, 249.994, 
    249.9938, 249.9942, 249.9939, 249.9944, 249.9935, 249.9939, 249.9931, 
    249.9932, 249.9934, 249.9937, 249.9935, 249.9937, 249.9933, 249.993, 
    249.993, 249.9928, 249.993, 249.993, 249.9931, 249.993, 249.9933, 
    249.9932, 249.9936, 249.9937, 249.9941, 249.9944, 249.9947, 249.9948, 
    249.9948, 249.9948 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.6145, 258.6148, 258.6148, 258.615, 258.6149, 258.6151, 258.6146, 
    258.6148, 258.6147, 258.6145, 258.6155, 258.615, 258.616, 258.6157, 
    258.6165, 258.616, 258.6166, 258.6165, 258.6168, 258.6167, 258.6172, 
    258.6169, 258.6174, 258.6171, 258.6171, 258.6169, 258.6151, 258.6154, 
    258.6151, 258.6151, 258.6151, 258.6149, 258.6147, 258.6145, 258.6145, 
    258.6147, 258.6152, 258.615, 258.6154, 258.6154, 258.6158, 258.6156, 
    258.6163, 258.6161, 258.6167, 258.6166, 258.6167, 258.6167, 258.6167, 
    258.6165, 258.6166, 258.6164, 258.6157, 258.6159, 258.6152, 258.6148, 
    258.6146, 258.6144, 258.6144, 258.6145, 258.6147, 258.615, 258.6151, 
    258.6153, 258.6154, 258.6158, 258.6159, 258.6164, 258.6163, 258.6164, 
    258.6165, 258.6168, 258.6167, 258.6168, 258.6164, 258.6167, 258.6163, 
    258.6164, 258.6154, 258.6151, 258.6149, 258.6148, 258.6144, 258.6147, 
    258.6146, 258.6148, 258.6149, 258.6149, 258.6153, 258.6151, 258.616, 
    258.6156, 258.6165, 258.6163, 258.6166, 258.6165, 258.6167, 258.6165, 
    258.6169, 258.6169, 258.6169, 258.6171, 258.6165, 258.6167, 258.6149, 
    258.6149, 258.6149, 258.6147, 258.6147, 258.6145, 258.6147, 258.6147, 
    258.615, 258.6151, 258.6152, 258.6154, 258.6157, 258.6161, 258.6163, 
    258.6165, 258.6164, 258.6165, 258.6164, 258.6163, 258.6169, 258.6166, 
    258.6171, 258.6171, 258.6168, 258.6171, 258.6149, 258.6148, 258.6146, 
    258.6148, 258.6145, 258.6147, 258.6147, 258.6151, 258.6152, 258.6153, 
    258.6154, 258.6156, 258.616, 258.6163, 258.6166, 258.6165, 258.6165, 
    258.6166, 258.6165, 258.6166, 258.6167, 258.6166, 258.617, 258.6169, 
    258.617, 258.617, 258.6148, 258.615, 258.6149, 258.615, 258.6149, 
    258.6153, 258.6154, 258.6158, 258.6156, 258.6159, 258.6157, 258.6157, 
    258.6159, 258.6157, 258.6163, 258.6159, 258.6166, 258.6162, 258.6166, 
    258.6166, 258.6167, 258.6168, 258.6169, 258.6172, 258.6172, 258.6174, 
    258.6151, 258.6152, 258.6152, 258.6154, 258.6155, 258.6157, 258.6161, 
    258.6159, 258.6162, 258.6162, 258.6158, 258.6161, 258.6153, 258.6154, 
    258.6154, 258.6151, 258.616, 258.6155, 258.6163, 258.6161, 258.6168, 
    258.6165, 258.6171, 258.6174, 258.6177, 258.618, 258.6153, 258.6152, 
    258.6154, 258.6156, 258.6158, 258.6161, 258.6161, 258.6162, 258.6163, 
    258.6165, 258.6162, 258.6165, 258.6155, 258.616, 258.6152, 258.6154, 
    258.6156, 258.6155, 258.6159, 258.616, 258.6164, 258.6162, 258.6173, 
    258.6168, 258.6183, 258.6179, 258.6152, 258.6153, 258.6158, 258.6155, 
    258.6161, 258.6163, 258.6164, 258.6165, 258.6166, 258.6166, 258.6165, 
    258.6166, 258.6161, 258.6164, 258.6157, 258.6158, 258.6158, 258.6157, 
    258.616, 258.6162, 258.6162, 258.6163, 258.6165, 258.6161, 258.6174, 
    258.6166, 258.6154, 258.6157, 258.6157, 258.6156, 258.6163, 258.616, 
    258.6166, 258.6165, 258.6168, 258.6166, 258.6166, 258.6164, 258.6163, 
    258.616, 258.6158, 258.6157, 258.6157, 258.6159, 258.6162, 258.6166, 
    258.6165, 258.6167, 258.6161, 258.6164, 258.6162, 258.6165, 258.6159, 
    258.6164, 258.6158, 258.6158, 258.616, 258.6164, 258.6165, 258.6165, 
    258.6165, 258.6162, 258.6162, 258.616, 258.616, 258.6158, 258.6157, 
    258.6158, 258.6159, 258.6162, 258.6165, 258.6168, 258.6169, 258.6172, 
    258.6169, 258.6174, 258.617, 258.6177, 258.6165, 258.617, 258.616, 
    258.6161, 258.6163, 258.6168, 258.6165, 258.6168, 258.6162, 258.6159, 
    258.6158, 258.6157, 258.6158, 258.6158, 258.6159, 258.6159, 258.6162, 
    258.6161, 258.6166, 258.6168, 258.6173, 258.6177, 258.618, 258.6182, 
    258.6183, 258.6183 ;

 TREFMXAV_R =
  258.6145, 258.6148, 258.6148, 258.615, 258.6149, 258.6151, 258.6146, 
    258.6148, 258.6147, 258.6145, 258.6155, 258.615, 258.616, 258.6157, 
    258.6165, 258.616, 258.6166, 258.6165, 258.6168, 258.6167, 258.6172, 
    258.6169, 258.6174, 258.6171, 258.6171, 258.6169, 258.6151, 258.6154, 
    258.6151, 258.6151, 258.6151, 258.6149, 258.6147, 258.6145, 258.6145, 
    258.6147, 258.6152, 258.615, 258.6154, 258.6154, 258.6158, 258.6156, 
    258.6163, 258.6161, 258.6167, 258.6166, 258.6167, 258.6167, 258.6167, 
    258.6165, 258.6166, 258.6164, 258.6157, 258.6159, 258.6152, 258.6148, 
    258.6146, 258.6144, 258.6144, 258.6145, 258.6147, 258.615, 258.6151, 
    258.6153, 258.6154, 258.6158, 258.6159, 258.6164, 258.6163, 258.6164, 
    258.6165, 258.6168, 258.6167, 258.6168, 258.6164, 258.6167, 258.6163, 
    258.6164, 258.6154, 258.6151, 258.6149, 258.6148, 258.6144, 258.6147, 
    258.6146, 258.6148, 258.6149, 258.6149, 258.6153, 258.6151, 258.616, 
    258.6156, 258.6165, 258.6163, 258.6166, 258.6165, 258.6167, 258.6165, 
    258.6169, 258.6169, 258.6169, 258.6171, 258.6165, 258.6167, 258.6149, 
    258.6149, 258.6149, 258.6147, 258.6147, 258.6145, 258.6147, 258.6147, 
    258.615, 258.6151, 258.6152, 258.6154, 258.6157, 258.6161, 258.6163, 
    258.6165, 258.6164, 258.6165, 258.6164, 258.6163, 258.6169, 258.6166, 
    258.6171, 258.6171, 258.6168, 258.6171, 258.6149, 258.6148, 258.6146, 
    258.6148, 258.6145, 258.6147, 258.6147, 258.6151, 258.6152, 258.6153, 
    258.6154, 258.6156, 258.616, 258.6163, 258.6166, 258.6165, 258.6165, 
    258.6166, 258.6165, 258.6166, 258.6167, 258.6166, 258.617, 258.6169, 
    258.617, 258.617, 258.6148, 258.615, 258.6149, 258.615, 258.6149, 
    258.6153, 258.6154, 258.6158, 258.6156, 258.6159, 258.6157, 258.6157, 
    258.6159, 258.6157, 258.6163, 258.6159, 258.6166, 258.6162, 258.6166, 
    258.6166, 258.6167, 258.6168, 258.6169, 258.6172, 258.6172, 258.6174, 
    258.6151, 258.6152, 258.6152, 258.6154, 258.6155, 258.6157, 258.6161, 
    258.6159, 258.6162, 258.6162, 258.6158, 258.6161, 258.6153, 258.6154, 
    258.6154, 258.6151, 258.616, 258.6155, 258.6163, 258.6161, 258.6168, 
    258.6165, 258.6171, 258.6174, 258.6177, 258.618, 258.6153, 258.6152, 
    258.6154, 258.6156, 258.6158, 258.6161, 258.6161, 258.6162, 258.6163, 
    258.6165, 258.6162, 258.6165, 258.6155, 258.616, 258.6152, 258.6154, 
    258.6156, 258.6155, 258.6159, 258.616, 258.6164, 258.6162, 258.6173, 
    258.6168, 258.6183, 258.6179, 258.6152, 258.6153, 258.6158, 258.6155, 
    258.6161, 258.6163, 258.6164, 258.6165, 258.6166, 258.6166, 258.6165, 
    258.6166, 258.6161, 258.6164, 258.6157, 258.6158, 258.6158, 258.6157, 
    258.616, 258.6162, 258.6162, 258.6163, 258.6165, 258.6161, 258.6174, 
    258.6166, 258.6154, 258.6157, 258.6157, 258.6156, 258.6163, 258.616, 
    258.6166, 258.6165, 258.6168, 258.6166, 258.6166, 258.6164, 258.6163, 
    258.616, 258.6158, 258.6157, 258.6157, 258.6159, 258.6162, 258.6166, 
    258.6165, 258.6167, 258.6161, 258.6164, 258.6162, 258.6165, 258.6159, 
    258.6164, 258.6158, 258.6158, 258.616, 258.6164, 258.6165, 258.6165, 
    258.6165, 258.6162, 258.6162, 258.616, 258.616, 258.6158, 258.6157, 
    258.6158, 258.6159, 258.6162, 258.6165, 258.6168, 258.6169, 258.6172, 
    258.6169, 258.6174, 258.617, 258.6177, 258.6165, 258.617, 258.616, 
    258.6161, 258.6163, 258.6168, 258.6165, 258.6168, 258.6162, 258.6159, 
    258.6158, 258.6157, 258.6158, 258.6158, 258.6159, 258.6159, 258.6162, 
    258.6161, 258.6166, 258.6168, 258.6173, 258.6177, 258.618, 258.6182, 
    258.6183, 258.6183 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.9799, 253.9801, 253.9801, 253.9802, 253.9801, 253.9802, 253.98, 
    253.9801, 253.98, 253.9799, 253.9804, 253.9802, 253.9807, 253.9805, 
    253.9809, 253.9807, 253.981, 253.9809, 253.9811, 253.981, 253.9813, 
    253.9811, 253.9814, 253.9812, 253.9813, 253.9811, 253.9802, 253.9804, 
    253.9802, 253.9803, 253.9802, 253.9801, 253.98, 253.9799, 253.9799, 
    253.98, 253.9803, 253.9802, 253.9804, 253.9804, 253.9806, 253.9805, 
    253.9809, 253.9808, 253.981, 253.981, 253.981, 253.981, 253.981, 
    253.9809, 253.981, 253.9809, 253.9805, 253.9806, 253.9803, 253.9801, 
    253.98, 253.9799, 253.9799, 253.9799, 253.98, 253.9802, 253.9803, 
    253.9803, 253.9804, 253.9805, 253.9807, 253.9809, 253.9808, 253.9809, 
    253.981, 253.9811, 253.9811, 253.9811, 253.9809, 253.981, 253.9808, 
    253.9809, 253.9804, 253.9802, 253.9801, 253.9801, 253.9799, 253.98, 
    253.98, 253.9801, 253.9801, 253.9801, 253.9803, 253.9802, 253.9807, 
    253.9805, 253.981, 253.9809, 253.981, 253.9809, 253.981, 253.9809, 
    253.9811, 253.9812, 253.9811, 253.9812, 253.9809, 253.981, 253.9801, 
    253.9801, 253.9801, 253.98, 253.98, 253.9799, 253.98, 253.98, 253.9801, 
    253.9802, 253.9803, 253.9804, 253.9805, 253.9807, 253.9809, 253.9809, 
    253.9809, 253.9809, 253.9809, 253.9809, 253.9811, 253.981, 253.9812, 
    253.9812, 253.9811, 253.9812, 253.9801, 253.9801, 253.98, 253.9801, 
    253.9799, 253.98, 253.98, 253.9802, 253.9803, 253.9803, 253.9804, 
    253.9805, 253.9807, 253.9808, 253.981, 253.981, 253.981, 253.981, 
    253.9809, 253.981, 253.981, 253.981, 253.9812, 253.9812, 253.9812, 
    253.9812, 253.9801, 253.9801, 253.9801, 253.9802, 253.9801, 253.9803, 
    253.9803, 253.9806, 253.9805, 253.9807, 253.9805, 253.9805, 253.9807, 
    253.9805, 253.9808, 253.9806, 253.981, 253.9808, 253.981, 253.981, 
    253.981, 253.9811, 253.9812, 253.9813, 253.9813, 253.9814, 253.9802, 
    253.9803, 253.9803, 253.9804, 253.9804, 253.9805, 253.9807, 253.9807, 
    253.9808, 253.9808, 253.9806, 253.9807, 253.9803, 253.9804, 253.9804, 
    253.9802, 253.9807, 253.9804, 253.9809, 253.9807, 253.9811, 253.9809, 
    253.9812, 253.9814, 253.9815, 253.9817, 253.9803, 253.9803, 253.9804, 
    253.9805, 253.9806, 253.9807, 253.9808, 253.9808, 253.9809, 253.9809, 
    253.9808, 253.9809, 253.9804, 253.9807, 253.9803, 253.9804, 253.9805, 
    253.9804, 253.9806, 253.9807, 253.9809, 253.9808, 253.9814, 253.9811, 
    253.9818, 253.9816, 253.9803, 253.9803, 253.9805, 253.9805, 253.9807, 
    253.9808, 253.9809, 253.981, 253.981, 253.981, 253.9809, 253.981, 
    253.9807, 253.9809, 253.9805, 253.9806, 253.9806, 253.9805, 253.9807, 
    253.9808, 253.9808, 253.9808, 253.9809, 253.9808, 253.9814, 253.981, 
    253.9804, 253.9805, 253.9805, 253.9805, 253.9808, 253.9807, 253.981, 
    253.9809, 253.9811, 253.981, 253.981, 253.9809, 253.9809, 253.9807, 
    253.9806, 253.9805, 253.9805, 253.9806, 253.9808, 253.981, 253.9809, 
    253.9811, 253.9807, 253.9809, 253.9808, 253.981, 253.9807, 253.9809, 
    253.9806, 253.9806, 253.9807, 253.9809, 253.9809, 253.981, 253.9809, 
    253.9808, 253.9808, 253.9807, 253.9807, 253.9806, 253.9805, 253.9806, 
    253.9807, 253.9808, 253.9809, 253.9811, 253.9811, 253.9813, 253.9812, 
    253.9814, 253.9812, 253.9815, 253.9809, 253.9812, 253.9807, 253.9808, 
    253.9809, 253.9811, 253.981, 253.9811, 253.9808, 253.9806, 253.9806, 
    253.9805, 253.9806, 253.9806, 253.9807, 253.9806, 253.9808, 253.9807, 
    253.981, 253.9811, 253.9814, 253.9815, 253.9817, 253.9818, 253.9818, 
    253.9818 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.9799, 253.9801, 253.9801, 253.9802, 253.9801, 253.9802, 253.98, 
    253.9801, 253.98, 253.9799, 253.9804, 253.9802, 253.9807, 253.9805, 
    253.9809, 253.9807, 253.981, 253.9809, 253.9811, 253.981, 253.9813, 
    253.9811, 253.9814, 253.9812, 253.9813, 253.9811, 253.9802, 253.9804, 
    253.9802, 253.9803, 253.9802, 253.9801, 253.98, 253.9799, 253.9799, 
    253.98, 253.9803, 253.9802, 253.9804, 253.9804, 253.9806, 253.9805, 
    253.9809, 253.9808, 253.981, 253.981, 253.981, 253.981, 253.981, 
    253.9809, 253.981, 253.9809, 253.9805, 253.9806, 253.9803, 253.9801, 
    253.98, 253.9799, 253.9799, 253.9799, 253.98, 253.9802, 253.9803, 
    253.9803, 253.9804, 253.9805, 253.9807, 253.9809, 253.9808, 253.9809, 
    253.981, 253.9811, 253.9811, 253.9811, 253.9809, 253.981, 253.9808, 
    253.9809, 253.9804, 253.9802, 253.9801, 253.9801, 253.9799, 253.98, 
    253.98, 253.9801, 253.9801, 253.9801, 253.9803, 253.9802, 253.9807, 
    253.9805, 253.981, 253.9809, 253.981, 253.9809, 253.981, 253.9809, 
    253.9811, 253.9812, 253.9811, 253.9812, 253.9809, 253.981, 253.9801, 
    253.9801, 253.9801, 253.98, 253.98, 253.9799, 253.98, 253.98, 253.9801, 
    253.9802, 253.9803, 253.9804, 253.9805, 253.9807, 253.9809, 253.9809, 
    253.9809, 253.9809, 253.9809, 253.9809, 253.9811, 253.981, 253.9812, 
    253.9812, 253.9811, 253.9812, 253.9801, 253.9801, 253.98, 253.9801, 
    253.9799, 253.98, 253.98, 253.9802, 253.9803, 253.9803, 253.9804, 
    253.9805, 253.9807, 253.9808, 253.981, 253.981, 253.981, 253.981, 
    253.9809, 253.981, 253.981, 253.981, 253.9812, 253.9812, 253.9812, 
    253.9812, 253.9801, 253.9801, 253.9801, 253.9802, 253.9801, 253.9803, 
    253.9803, 253.9806, 253.9805, 253.9807, 253.9805, 253.9805, 253.9807, 
    253.9805, 253.9808, 253.9806, 253.981, 253.9808, 253.981, 253.981, 
    253.981, 253.9811, 253.9812, 253.9813, 253.9813, 253.9814, 253.9802, 
    253.9803, 253.9803, 253.9804, 253.9804, 253.9805, 253.9807, 253.9807, 
    253.9808, 253.9808, 253.9806, 253.9807, 253.9803, 253.9804, 253.9804, 
    253.9802, 253.9807, 253.9804, 253.9809, 253.9807, 253.9811, 253.9809, 
    253.9812, 253.9814, 253.9815, 253.9817, 253.9803, 253.9803, 253.9804, 
    253.9805, 253.9806, 253.9807, 253.9808, 253.9808, 253.9809, 253.9809, 
    253.9808, 253.9809, 253.9804, 253.9807, 253.9803, 253.9804, 253.9805, 
    253.9804, 253.9806, 253.9807, 253.9809, 253.9808, 253.9814, 253.9811, 
    253.9818, 253.9816, 253.9803, 253.9803, 253.9805, 253.9805, 253.9807, 
    253.9808, 253.9809, 253.981, 253.981, 253.981, 253.9809, 253.981, 
    253.9807, 253.9809, 253.9805, 253.9806, 253.9806, 253.9805, 253.9807, 
    253.9808, 253.9808, 253.9808, 253.9809, 253.9808, 253.9814, 253.981, 
    253.9804, 253.9805, 253.9805, 253.9805, 253.9808, 253.9807, 253.981, 
    253.9809, 253.9811, 253.981, 253.981, 253.9809, 253.9809, 253.9807, 
    253.9806, 253.9805, 253.9805, 253.9806, 253.9808, 253.981, 253.9809, 
    253.9811, 253.9807, 253.9809, 253.9808, 253.981, 253.9807, 253.9809, 
    253.9806, 253.9806, 253.9807, 253.9809, 253.9809, 253.981, 253.9809, 
    253.9808, 253.9808, 253.9807, 253.9807, 253.9806, 253.9805, 253.9806, 
    253.9807, 253.9808, 253.9809, 253.9811, 253.9811, 253.9813, 253.9812, 
    253.9814, 253.9812, 253.9815, 253.9809, 253.9812, 253.9807, 253.9808, 
    253.9809, 253.9811, 253.981, 253.9811, 253.9808, 253.9806, 253.9806, 
    253.9805, 253.9806, 253.9806, 253.9807, 253.9806, 253.9808, 253.9807, 
    253.981, 253.9811, 253.9814, 253.9815, 253.9817, 253.9818, 253.9818, 
    253.9818 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.5822, 254.5837, 254.5834, 254.5846, 254.584, 254.5847, 254.5825, 
    254.5837, 254.583, 254.5824, 254.5868, 254.5847, 254.5892, 254.5878, 
    254.5914, 254.589, 254.5919, 254.5914, 254.5931, 254.5926, 254.5947, 
    254.5933, 254.5959, 254.5944, 254.5946, 254.5933, 254.5851, 254.5865, 
    254.585, 254.5852, 254.5851, 254.584, 254.5833, 254.5821, 254.5824, 
    254.5833, 254.5853, 254.5846, 254.5864, 254.5864, 254.5884, 254.5875, 
    254.5908, 254.5899, 254.5927, 254.5919, 254.5926, 254.5924, 254.5926, 
    254.5916, 254.592, 254.5911, 254.5876, 254.5887, 254.5856, 254.5837, 
    254.5826, 254.5817, 254.5818, 254.5821, 254.5833, 254.5844, 254.5853, 
    254.5858, 254.5864, 254.588, 254.589, 254.591, 254.5907, 254.5913, 
    254.5919, 254.5929, 254.5927, 254.5931, 254.5913, 254.5925, 254.5905, 
    254.591, 254.5864, 254.5848, 254.5841, 254.5835, 254.5819, 254.583, 
    254.5826, 254.5836, 254.5842, 254.5839, 254.5858, 254.5851, 254.589, 
    254.5873, 254.5918, 254.5907, 254.5921, 254.5914, 254.5925, 254.5915, 
    254.5933, 254.5937, 254.5934, 254.5945, 254.5914, 254.5926, 254.5839, 
    254.5839, 254.5842, 254.5831, 254.5831, 254.5821, 254.583, 254.5833, 
    254.5843, 254.5848, 254.5853, 254.5865, 254.5877, 254.5895, 254.5908, 
    254.5917, 254.5911, 254.5916, 254.5911, 254.5909, 254.5935, 254.592, 
    254.5943, 254.5942, 254.5932, 254.5942, 254.584, 254.5837, 254.5827, 
    254.5835, 254.582, 254.5828, 254.5833, 254.5851, 254.5855, 254.5859, 
    254.5866, 254.5875, 254.5892, 254.5906, 254.5919, 254.5918, 254.5919, 
    254.5921, 254.5914, 254.5923, 254.5924, 254.592, 254.5942, 254.5936, 
    254.5942, 254.5938, 254.5838, 254.5843, 254.584, 254.5845, 254.5842, 
    254.5857, 254.5862, 254.5884, 254.5875, 254.5889, 254.5876, 254.5879, 
    254.5889, 254.5877, 254.5905, 254.5886, 254.5921, 254.5902, 254.5923, 
    254.5919, 254.5925, 254.593, 254.5938, 254.595, 254.5947, 254.5958, 
    254.585, 254.5856, 254.5856, 254.5863, 254.5868, 254.5878, 254.5896, 
    254.5889, 254.5901, 254.5904, 254.5885, 254.5896, 254.5861, 254.5866, 
    254.5863, 254.5851, 254.5891, 254.587, 254.5908, 254.5897, 254.593, 
    254.5913, 254.5945, 254.5959, 254.5972, 254.5987, 254.586, 254.5856, 
    254.5863, 254.5874, 254.5884, 254.5898, 254.5899, 254.5902, 254.5908, 
    254.5914, 254.5902, 254.5915, 254.5867, 254.5892, 254.5854, 254.5865, 
    254.5873, 254.587, 254.5889, 254.5893, 254.591, 254.5901, 254.5955, 
    254.5931, 254.5999, 254.598, 254.5854, 254.586, 254.588, 254.5871, 
    254.5899, 254.5905, 254.5911, 254.5918, 254.5919, 254.5923, 254.5916, 
    254.5923, 254.5898, 254.5909, 254.5878, 254.5886, 254.5882, 254.5878, 
    254.589, 254.5902, 254.5903, 254.5907, 254.5917, 254.5899, 254.5958, 
    254.5921, 254.5867, 254.5877, 254.5879, 254.5875, 254.5905, 254.5894, 
    254.5923, 254.5915, 254.5928, 254.5922, 254.5921, 254.5913, 254.5907, 
    254.5894, 254.5884, 254.5876, 254.5878, 254.5887, 254.5903, 254.5919, 
    254.5916, 254.5927, 254.5897, 254.5909, 254.5904, 254.5917, 254.5889, 
    254.5912, 254.5883, 254.5886, 254.5894, 254.591, 254.5914, 254.5918, 
    254.5916, 254.5904, 254.5902, 254.5894, 254.5891, 254.5885, 254.588, 
    254.5885, 254.5889, 254.5904, 254.5916, 254.593, 254.5934, 254.595, 
    254.5937, 254.5958, 254.5939, 254.5972, 254.5914, 254.5939, 254.5894, 
    254.5899, 254.5908, 254.5928, 254.5917, 254.593, 254.5902, 254.5887, 
    254.5883, 254.5876, 254.5883, 254.5883, 254.589, 254.5888, 254.5904, 
    254.5895, 254.5921, 254.593, 254.5956, 254.5972, 254.5989, 254.5997, 
    254.5999, 254.6,
  255.7167, 255.7182, 255.7179, 255.7192, 255.7185, 255.7193, 255.717, 
    255.7183, 255.7175, 255.7169, 255.7215, 255.7192, 255.724, 255.7225, 
    255.7263, 255.7238, 255.7269, 255.7263, 255.7281, 255.7276, 255.7298, 
    255.7283, 255.731, 255.7294, 255.7297, 255.7282, 255.7197, 255.7212, 
    255.7196, 255.7198, 255.7197, 255.7185, 255.7179, 255.7166, 255.7168, 
    255.7178, 255.7199, 255.7192, 255.7211, 255.7211, 255.7231, 255.7222, 
    255.7257, 255.7247, 255.7276, 255.7269, 255.7275, 255.7273, 255.7275, 
    255.7265, 255.7269, 255.726, 255.7224, 255.7234, 255.7202, 255.7183, 
    255.7171, 255.7162, 255.7163, 255.7166, 255.7178, 255.719, 255.7198, 
    255.7204, 255.721, 255.7227, 255.7237, 255.7259, 255.7255, 255.7261, 
    255.7268, 255.7278, 255.7276, 255.7281, 255.7261, 255.7274, 255.7253, 
    255.7259, 255.7211, 255.7194, 255.7186, 255.718, 255.7164, 255.7175, 
    255.7171, 255.7181, 255.7188, 255.7185, 255.7205, 255.7197, 255.7238, 
    255.722, 255.7267, 255.7256, 255.727, 255.7263, 255.7275, 255.7264, 
    255.7283, 255.7287, 255.7284, 255.7295, 255.7263, 255.7275, 255.7184, 
    255.7185, 255.7187, 255.7176, 255.7176, 255.7166, 255.7175, 255.7178, 
    255.7188, 255.7194, 255.7199, 255.7211, 255.7224, 255.7243, 255.7256, 
    255.7266, 255.726, 255.7265, 255.726, 255.7257, 255.7285, 255.7269, 
    255.7293, 255.7292, 255.7281, 255.7292, 255.7185, 255.7182, 255.7172, 
    255.718, 255.7165, 255.7173, 255.7178, 255.7197, 255.7201, 255.7205, 
    255.7213, 255.7222, 255.7239, 255.7254, 255.7268, 255.7267, 255.7267, 
    255.7271, 255.7263, 255.7272, 255.7273, 255.7269, 255.7292, 255.7285, 
    255.7292, 255.7288, 255.7183, 255.7188, 255.7186, 255.7191, 255.7187, 
    255.7203, 255.7208, 255.7231, 255.7222, 255.7237, 255.7224, 255.7226, 
    255.7237, 255.7224, 255.7253, 255.7233, 255.7271, 255.725, 255.7272, 
    255.7268, 255.7274, 255.728, 255.7287, 255.73, 255.7297, 255.7309, 
    255.7196, 255.7203, 255.7202, 255.7209, 255.7214, 255.7226, 255.7244, 
    255.7237, 255.7249, 255.7252, 255.7233, 255.7244, 255.7207, 255.7213, 
    255.721, 255.7197, 255.7238, 255.7217, 255.7257, 255.7245, 255.7279, 
    255.7262, 255.7296, 255.731, 255.7324, 255.7339, 255.7206, 255.7202, 
    255.721, 255.7221, 255.7232, 255.7246, 255.7247, 255.725, 255.7257, 
    255.7262, 255.725, 255.7264, 255.7214, 255.724, 255.72, 255.7212, 
    255.722, 255.7217, 255.7236, 255.7241, 255.7259, 255.725, 255.7306, 
    255.7281, 255.7352, 255.7332, 255.72, 255.7206, 255.7227, 255.7218, 
    255.7247, 255.7254, 255.726, 255.7267, 255.7268, 255.7272, 255.7265, 
    255.7272, 255.7246, 255.7258, 255.7225, 255.7233, 255.723, 255.7226, 
    255.7238, 255.7251, 255.7251, 255.7255, 255.7266, 255.7247, 255.7309, 
    255.727, 255.7213, 255.7225, 255.7227, 255.7222, 255.7253, 255.7242, 
    255.7272, 255.7264, 255.7278, 255.7271, 255.727, 255.7261, 255.7256, 
    255.7242, 255.7231, 255.7223, 255.7225, 255.7234, 255.7251, 255.7268, 
    255.7264, 255.7277, 255.7245, 255.7258, 255.7253, 255.7266, 255.7237, 
    255.7261, 255.723, 255.7233, 255.7242, 255.7259, 255.7263, 255.7267, 
    255.7264, 255.7252, 255.725, 255.7242, 255.7239, 255.7233, 255.7227, 
    255.7232, 255.7237, 255.7252, 255.7265, 255.728, 255.7284, 255.73, 
    255.7287, 255.7309, 255.7289, 255.7324, 255.7263, 255.7289, 255.7242, 
    255.7247, 255.7256, 255.7278, 255.7266, 255.728, 255.725, 255.7234, 
    255.7231, 255.7223, 255.7231, 255.723, 255.7238, 255.7235, 255.7253, 
    255.7243, 255.727, 255.728, 255.7307, 255.7324, 255.7342, 255.735, 
    255.7352, 255.7353,
  257.2881, 257.2897, 257.2894, 257.2907, 257.29, 257.2909, 257.2884, 
    257.2898, 257.2889, 257.2882, 257.2933, 257.2908, 257.2961, 257.2944, 
    257.2986, 257.2958, 257.2991, 257.2985, 257.3004, 257.2999, 257.3023, 
    257.3007, 257.3036, 257.3019, 257.3022, 257.3006, 257.2914, 257.293, 
    257.2912, 257.2915, 257.2914, 257.29, 257.2893, 257.288, 257.2882, 
    257.2892, 257.2916, 257.2908, 257.2928, 257.2928, 257.295, 257.294, 
    257.2978, 257.2968, 257.2999, 257.2991, 257.2999, 257.2996, 257.2999, 
    257.2987, 257.2992, 257.2982, 257.2942, 257.2953, 257.2919, 257.2898, 
    257.2885, 257.2875, 257.2876, 257.2879, 257.2892, 257.2905, 257.2915, 
    257.2921, 257.2928, 257.2946, 257.2957, 257.298, 257.2976, 257.2983, 
    257.299, 257.3002, 257.3, 257.3005, 257.2983, 257.2997, 257.2974, 
    257.298, 257.2929, 257.291, 257.2902, 257.2895, 257.2878, 257.2889, 
    257.2885, 257.2896, 257.2903, 257.2899, 257.2921, 257.2913, 257.2958, 
    257.2939, 257.299, 257.2977, 257.2993, 257.2985, 257.2998, 257.2986, 
    257.3007, 257.3011, 257.3008, 257.302, 257.2985, 257.2999, 257.2899, 
    257.29, 257.2903, 257.2891, 257.289, 257.2879, 257.2889, 257.2893, 
    257.2903, 257.291, 257.2916, 257.2928, 257.2943, 257.2963, 257.2978, 
    257.2988, 257.2982, 257.2987, 257.2981, 257.2979, 257.3009, 257.2992, 
    257.3018, 257.3017, 257.3005, 257.3017, 257.29, 257.2897, 257.2885, 
    257.2895, 257.2878, 257.2887, 257.2892, 257.2913, 257.2918, 257.2922, 
    257.293, 257.2941, 257.2959, 257.2975, 257.2991, 257.299, 257.299, 
    257.2993, 257.2985, 257.2995, 257.2996, 257.2992, 257.3017, 257.301, 
    257.3017, 257.3012, 257.2898, 257.2904, 257.2901, 257.2906, 257.2903, 
    257.292, 257.2925, 257.295, 257.294, 257.2957, 257.2942, 257.2945, 
    257.2957, 257.2943, 257.2975, 257.2953, 257.2993, 257.2971, 257.2995, 
    257.2991, 257.2997, 257.3004, 257.3011, 257.3026, 257.3023, 257.3035, 
    257.2912, 257.2919, 257.2919, 257.2926, 257.2932, 257.2944, 257.2964, 
    257.2957, 257.297, 257.2973, 257.2952, 257.2965, 257.2924, 257.2931, 
    257.2927, 257.2913, 257.2958, 257.2935, 257.2978, 257.2965, 257.3003, 
    257.2984, 257.3021, 257.3036, 257.3051, 257.3068, 257.2923, 257.2918, 
    257.2927, 257.2939, 257.2951, 257.2966, 257.2968, 257.2971, 257.2978, 
    257.2984, 257.2971, 257.2986, 257.2932, 257.296, 257.2917, 257.2929, 
    257.2939, 257.2935, 257.2956, 257.2961, 257.2981, 257.2971, 257.3032, 
    257.3005, 257.3082, 257.306, 257.2917, 257.2924, 257.2946, 257.2935, 
    257.2967, 257.2975, 257.2982, 257.299, 257.2991, 257.2995, 257.2988, 
    257.2995, 257.2966, 257.2979, 257.2944, 257.2953, 257.2949, 257.2944, 
    257.2958, 257.2971, 257.2972, 257.2977, 257.2989, 257.2968, 257.3035, 
    257.2993, 257.2931, 257.2943, 257.2945, 257.294, 257.2974, 257.2962, 
    257.2995, 257.2986, 257.3001, 257.2994, 257.2993, 257.2983, 257.2977, 
    257.2963, 257.295, 257.2941, 257.2943, 257.2954, 257.2972, 257.2991, 
    257.2986, 257.3, 257.2965, 257.2979, 257.2974, 257.2989, 257.2957, 
    257.2983, 257.295, 257.2953, 257.2962, 257.298, 257.2985, 257.2989, 
    257.2986, 257.2973, 257.2971, 257.2962, 257.2959, 257.2952, 257.2946, 
    257.2951, 257.2957, 257.2973, 257.2988, 257.3004, 257.3008, 257.3026, 
    257.3011, 257.3035, 257.3014, 257.3051, 257.2985, 257.3014, 257.2962, 
    257.2968, 257.2978, 257.3001, 257.2989, 257.3003, 257.2971, 257.2954, 
    257.295, 257.2942, 257.295, 257.2949, 257.2957, 257.2955, 257.2974, 
    257.2964, 257.2993, 257.3003, 257.3033, 257.3052, 257.3071, 257.308, 
    257.3082, 257.3083,
  259.3232, 259.3249, 259.3246, 259.326, 259.3252, 259.3261, 259.3236, 
    259.325, 259.3241, 259.3234, 259.3286, 259.326, 259.3314, 259.3297, 
    259.3339, 259.3311, 259.3345, 259.3339, 259.3358, 259.3353, 259.3377, 
    259.3361, 259.3391, 259.3373, 259.3376, 259.336, 259.3266, 259.3283, 
    259.3264, 259.3267, 259.3266, 259.3252, 259.3245, 259.3231, 259.3234, 
    259.3244, 259.3268, 259.326, 259.3281, 259.328, 259.3303, 259.3293, 
    259.3332, 259.3321, 259.3353, 259.3345, 259.3352, 259.335, 259.3352, 
    259.334, 259.3346, 259.3335, 259.3295, 259.3307, 259.3271, 259.325, 
    259.3236, 259.3227, 259.3228, 259.3231, 259.3244, 259.3257, 259.3267, 
    259.3274, 259.328, 259.33, 259.331, 259.3334, 259.333, 259.3337, 
    259.3344, 259.3355, 259.3354, 259.3359, 259.3337, 259.3351, 259.3327, 
    259.3334, 259.3281, 259.3262, 259.3253, 259.3246, 259.3229, 259.3241, 
    259.3236, 259.3248, 259.3255, 259.3252, 259.3274, 259.3265, 259.3311, 
    259.3291, 259.3343, 259.3331, 259.3346, 259.3338, 259.3352, 259.334, 
    259.3361, 259.3365, 259.3362, 259.3374, 259.3339, 259.3352, 259.3251, 
    259.3252, 259.3255, 259.3242, 259.3242, 259.3231, 259.3241, 259.3245, 
    259.3256, 259.3262, 259.3268, 259.3281, 259.3296, 259.3316, 259.3331, 
    259.3341, 259.3335, 259.3341, 259.3335, 259.3332, 259.3363, 259.3346, 
    259.3372, 259.3371, 259.3359, 259.3371, 259.3252, 259.3249, 259.3237, 
    259.3246, 259.323, 259.3239, 259.3244, 259.3265, 259.327, 259.3274, 
    259.3282, 259.3293, 259.3312, 259.3329, 259.3344, 259.3343, 259.3344, 
    259.3347, 259.3339, 259.3348, 259.335, 259.3346, 259.3371, 259.3364, 
    259.3371, 259.3366, 259.325, 259.3256, 259.3253, 259.3258, 259.3254, 
    259.3272, 259.3278, 259.3304, 259.3293, 259.331, 259.3295, 259.3297, 
    259.331, 259.3296, 259.3328, 259.3306, 259.3347, 259.3325, 259.3348, 
    259.3344, 259.3351, 259.3358, 259.3365, 259.338, 259.3377, 259.3389, 
    259.3264, 259.3271, 259.3271, 259.3279, 259.3285, 259.3297, 259.3317, 
    259.331, 259.3323, 259.3326, 259.3305, 259.3318, 259.3277, 259.3283, 
    259.3279, 259.3265, 259.3311, 259.3287, 259.3332, 259.3318, 259.3357, 
    259.3338, 259.3375, 259.3391, 259.3406, 259.3424, 259.3276, 259.3271, 
    259.328, 259.3292, 259.3304, 259.3319, 259.3321, 259.3324, 259.3332, 
    259.3338, 259.3325, 259.334, 259.3284, 259.3313, 259.3269, 259.3282, 
    259.3291, 259.3287, 259.3309, 259.3314, 259.3334, 259.3324, 259.3387, 
    259.3359, 259.3438, 259.3415, 259.3269, 259.3276, 259.3299, 259.3288, 
    259.332, 259.3328, 259.3335, 259.3343, 259.3344, 259.3349, 259.3341, 
    259.3349, 259.3319, 259.3333, 259.3297, 259.3305, 259.3301, 259.3297, 
    259.3311, 259.3325, 259.3326, 259.333, 259.3343, 259.3321, 259.339, 
    259.3347, 259.3283, 259.3296, 259.3298, 259.3293, 259.3328, 259.3315, 
    259.3349, 259.334, 259.3355, 259.3347, 259.3346, 259.3337, 259.3331, 
    259.3315, 259.3303, 259.3294, 259.3296, 259.3307, 259.3326, 259.3344, 
    259.334, 259.3354, 259.3318, 259.3333, 259.3327, 259.3342, 259.3309, 
    259.3337, 259.3302, 259.3305, 259.3315, 259.3334, 259.3338, 259.3343, 
    259.334, 259.3326, 259.3324, 259.3315, 259.3312, 259.3305, 259.3299, 
    259.3304, 259.331, 259.3326, 259.3341, 259.3358, 259.3362, 259.338, 
    259.3365, 259.339, 259.3368, 259.3407, 259.3339, 259.3368, 259.3315, 
    259.3321, 259.3331, 259.3355, 259.3342, 259.3357, 259.3324, 259.3307, 
    259.3303, 259.3294, 259.3303, 259.3302, 259.331, 259.3307, 259.3327, 
    259.3317, 259.3346, 259.3357, 259.3388, 259.3407, 259.3427, 259.3435, 
    259.3438, 259.3439,
  261.4319, 261.4331, 261.4329, 261.4339, 261.4333, 261.4341, 261.4321, 
    261.4332, 261.4325, 261.432, 261.436, 261.434, 261.4381, 261.4368, 
    261.4401, 261.4379, 261.4405, 261.44, 261.4415, 261.4411, 261.443, 
    261.4417, 261.444, 261.4427, 261.4429, 261.4417, 261.4344, 261.4357, 
    261.4343, 261.4345, 261.4344, 261.4334, 261.4328, 261.4318, 261.4319, 
    261.4327, 261.4346, 261.434, 261.4355, 261.4355, 261.4373, 261.4365, 
    261.4395, 261.4386, 261.4411, 261.4405, 261.4411, 261.4409, 261.4411, 
    261.4402, 261.4406, 261.4397, 261.4366, 261.4375, 261.4348, 261.4332, 
    261.4322, 261.4314, 261.4315, 261.4317, 261.4328, 261.4337, 261.4345, 
    261.435, 261.4355, 261.437, 261.4378, 261.4396, 261.4393, 261.4399, 
    261.4404, 261.4413, 261.4412, 261.4416, 261.4398, 261.441, 261.4391, 
    261.4396, 261.4356, 261.4341, 261.4335, 261.433, 261.4316, 261.4325, 
    261.4322, 261.433, 261.4336, 261.4333, 261.435, 261.4344, 261.4379, 
    261.4364, 261.4403, 261.4394, 261.4406, 261.44, 261.441, 261.4401, 
    261.4417, 261.442, 261.4418, 261.4427, 261.44, 261.4411, 261.4333, 
    261.4333, 261.4336, 261.4326, 261.4326, 261.4317, 261.4325, 261.4328, 
    261.4336, 261.4341, 261.4346, 261.4356, 261.4367, 261.4383, 261.4395, 
    261.4402, 261.4398, 261.4402, 261.4397, 261.4395, 261.4419, 261.4406, 
    261.4426, 261.4425, 261.4416, 261.4425, 261.4334, 261.4331, 261.4322, 
    261.4329, 261.4316, 261.4324, 261.4328, 261.4344, 261.4347, 261.4351, 
    261.4357, 261.4365, 261.438, 261.4393, 261.4404, 261.4403, 261.4404, 
    261.4406, 261.44, 261.4407, 261.4409, 261.4406, 261.4425, 261.4419, 
    261.4425, 261.4421, 261.4332, 261.4337, 261.4334, 261.4338, 261.4335, 
    261.4349, 261.4353, 261.4373, 261.4365, 261.4378, 261.4366, 261.4368, 
    261.4378, 261.4367, 261.4392, 261.4375, 261.4406, 261.4389, 261.4408, 
    261.4404, 261.441, 261.4415, 261.4421, 261.4432, 261.443, 261.4439, 
    261.4343, 261.4349, 261.4348, 261.4354, 261.4359, 261.4368, 261.4384, 
    261.4378, 261.4388, 261.4391, 261.4374, 261.4384, 261.4352, 261.4358, 
    261.4355, 261.4344, 261.4379, 261.4361, 261.4395, 261.4385, 261.4414, 
    261.4399, 261.4428, 261.444, 261.4452, 261.4466, 261.4352, 261.4348, 
    261.4355, 261.4364, 261.4373, 261.4385, 261.4387, 261.4389, 261.4395, 
    261.4399, 261.4389, 261.4401, 261.4359, 261.438, 261.4346, 261.4357, 
    261.4364, 261.4361, 261.4377, 261.4381, 261.4397, 261.4388, 261.4437, 
    261.4416, 261.4476, 261.4459, 261.4347, 261.4352, 261.437, 261.4361, 
    261.4386, 261.4392, 261.4397, 261.4404, 261.4404, 261.4408, 261.4402, 
    261.4408, 261.4385, 261.4395, 261.4368, 261.4374, 261.4371, 261.4368, 
    261.4379, 261.439, 261.439, 261.4393, 261.4403, 261.4386, 261.444, 
    261.4406, 261.4358, 261.4367, 261.4369, 261.4365, 261.4391, 261.4382, 
    261.4408, 261.4401, 261.4413, 261.4407, 261.4406, 261.4398, 261.4394, 
    261.4382, 261.4373, 261.4366, 261.4367, 261.4375, 261.439, 261.4404, 
    261.4401, 261.4412, 261.4384, 261.4396, 261.4391, 261.4403, 261.4377, 
    261.4399, 261.4372, 261.4374, 261.4382, 261.4396, 261.44, 261.4403, 
    261.4401, 261.4391, 261.4389, 261.4382, 261.438, 261.4374, 261.4369, 
    261.4373, 261.4378, 261.4391, 261.4402, 261.4415, 261.4418, 261.4432, 
    261.442, 261.444, 261.4423, 261.4453, 261.44, 261.4423, 261.4382, 
    261.4387, 261.4394, 261.4413, 261.4403, 261.4414, 261.4389, 261.4376, 
    261.4372, 261.4366, 261.4373, 261.4372, 261.4378, 261.4376, 261.4391, 
    261.4383, 261.4406, 261.4414, 261.4438, 261.4453, 261.4468, 261.4474, 
    261.4476, 261.4477,
  262.7628, 262.7633, 262.7632, 262.7636, 262.7634, 262.7637, 262.7629, 
    262.7633, 262.7631, 262.7629, 262.7645, 262.7637, 262.7653, 262.7648, 
    262.7661, 262.7652, 262.7662, 262.7661, 262.7666, 262.7664, 262.7672, 
    262.7667, 262.7676, 262.7671, 262.7672, 262.7667, 262.7638, 262.7643, 
    262.7638, 262.7639, 262.7638, 262.7634, 262.7632, 262.7628, 262.7628, 
    262.7632, 262.7639, 262.7637, 262.7643, 262.7643, 262.765, 262.7646, 
    262.7658, 262.7655, 262.7665, 262.7662, 262.7664, 262.7664, 262.7664, 
    262.7661, 262.7663, 262.7659, 262.7647, 262.7651, 262.764, 262.7634, 
    262.7629, 262.7626, 262.7627, 262.7628, 262.7632, 262.7636, 262.7639, 
    262.7641, 262.7643, 262.7649, 262.7652, 262.7659, 262.7658, 262.766, 
    262.7662, 262.7665, 262.7665, 262.7667, 262.766, 262.7664, 262.7657, 
    262.7659, 262.7643, 262.7637, 262.7635, 262.7632, 262.7627, 262.7631, 
    262.7629, 262.7633, 262.7635, 262.7634, 262.7641, 262.7638, 262.7652, 
    262.7646, 262.7662, 262.7658, 262.7663, 262.766, 262.7664, 262.7661, 
    262.7667, 262.7668, 262.7668, 262.7671, 262.7661, 262.7664, 262.7634, 
    262.7634, 262.7635, 262.7631, 262.7631, 262.7628, 262.7631, 262.7632, 
    262.7635, 262.7637, 262.7639, 262.7643, 262.7647, 262.7654, 262.7658, 
    262.7661, 262.7659, 262.7661, 262.7659, 262.7658, 262.7668, 262.7663, 
    262.7671, 262.767, 262.7667, 262.767, 262.7634, 262.7633, 262.763, 
    262.7632, 262.7628, 262.763, 262.7632, 262.7638, 262.7639, 262.7641, 
    262.7643, 262.7647, 262.7652, 262.7657, 262.7662, 262.7662, 262.7662, 
    262.7663, 262.766, 262.7663, 262.7664, 262.7663, 262.767, 262.7668, 
    262.767, 262.7669, 262.7634, 262.7635, 262.7634, 262.7636, 262.7635, 
    262.764, 262.7642, 262.765, 262.7646, 262.7652, 262.7647, 262.7648, 
    262.7652, 262.7647, 262.7657, 262.765, 262.7663, 262.7656, 262.7663, 
    262.7662, 262.7664, 262.7666, 262.7669, 262.7673, 262.7672, 262.7676, 
    262.7638, 262.764, 262.764, 262.7642, 262.7644, 262.7648, 262.7654, 
    262.7652, 262.7656, 262.7657, 262.765, 262.7654, 262.7642, 262.7644, 
    262.7643, 262.7638, 262.7652, 262.7645, 262.7658, 262.7654, 262.7666, 
    262.766, 262.7672, 262.7676, 262.7681, 262.7686, 262.7641, 262.764, 
    262.7643, 262.7646, 262.765, 262.7654, 262.7655, 262.7656, 262.7658, 
    262.766, 262.7656, 262.7661, 262.7644, 262.7653, 262.7639, 262.7643, 
    262.7646, 262.7645, 262.7651, 262.7653, 262.7659, 262.7656, 262.7675, 
    262.7667, 262.769, 262.7684, 262.7639, 262.7641, 262.7649, 262.7645, 
    262.7655, 262.7657, 262.7659, 262.7662, 262.7662, 262.7664, 262.7661, 
    262.7664, 262.7655, 262.7659, 262.7648, 262.765, 262.7649, 262.7648, 
    262.7652, 262.7656, 262.7656, 262.7658, 262.7662, 262.7655, 262.7676, 
    262.7663, 262.7643, 262.7647, 262.7648, 262.7646, 262.7657, 262.7653, 
    262.7664, 262.7661, 262.7665, 262.7663, 262.7663, 262.766, 262.7658, 
    262.7654, 262.765, 262.7647, 262.7647, 262.7651, 262.7657, 262.7662, 
    262.7661, 262.7665, 262.7654, 262.7659, 262.7657, 262.7661, 262.7652, 
    262.766, 262.7649, 262.765, 262.7653, 262.7659, 262.766, 262.7662, 
    262.7661, 262.7657, 262.7656, 262.7653, 262.7652, 262.765, 262.7648, 
    262.765, 262.7652, 262.7657, 262.7661, 262.7666, 262.7668, 262.7673, 
    262.7668, 262.7676, 262.767, 262.7681, 262.7661, 262.7669, 262.7653, 
    262.7655, 262.7658, 262.7665, 262.7661, 262.7666, 262.7656, 262.7651, 
    262.765, 262.7647, 262.765, 262.7649, 262.7652, 262.7651, 262.7657, 
    262.7654, 262.7663, 262.7666, 262.7675, 262.7681, 262.7687, 262.769, 
    262.7691, 262.7691,
  263.1171, 263.1172, 263.1171, 263.1172, 263.1172, 263.1172, 263.1171, 
    263.1172, 263.1171, 263.1171, 263.1173, 263.1172, 263.1174, 263.1174, 
    263.1176, 263.1174, 263.1176, 263.1176, 263.1176, 263.1176, 263.1177, 
    263.1176, 263.1178, 263.1177, 263.1177, 263.1176, 263.1172, 263.1173, 
    263.1172, 263.1172, 263.1172, 263.1172, 263.1171, 263.1171, 263.1171, 
    263.1171, 263.1172, 263.1172, 263.1173, 263.1173, 263.1174, 263.1173, 
    263.1175, 263.1175, 263.1176, 263.1176, 263.1176, 263.1176, 263.1176, 
    263.1176, 263.1176, 263.1176, 263.1174, 263.1174, 263.1172, 263.1172, 
    263.1171, 263.1171, 263.1171, 263.1171, 263.1171, 263.1172, 263.1172, 
    263.1172, 263.1173, 263.1174, 263.1174, 263.1175, 263.1175, 263.1176, 
    263.1176, 263.1176, 263.1176, 263.1176, 263.1176, 263.1176, 263.1175, 
    263.1175, 263.1173, 263.1172, 263.1172, 263.1172, 263.1171, 263.1171, 
    263.1171, 263.1172, 263.1172, 263.1172, 263.1173, 263.1172, 263.1174, 
    263.1173, 263.1176, 263.1175, 263.1176, 263.1176, 263.1176, 263.1176, 
    263.1176, 263.1177, 263.1176, 263.1177, 263.1176, 263.1176, 263.1172, 
    263.1172, 263.1172, 263.1171, 263.1171, 263.1171, 263.1171, 263.1171, 
    263.1172, 263.1172, 263.1172, 263.1173, 263.1174, 263.1175, 263.1175, 
    263.1176, 263.1176, 263.1176, 263.1175, 263.1175, 263.1177, 263.1176, 
    263.1177, 263.1177, 263.1176, 263.1177, 263.1172, 263.1172, 263.1171, 
    263.1172, 263.1171, 263.1171, 263.1171, 263.1172, 263.1172, 263.1173, 
    263.1173, 263.1173, 263.1174, 263.1175, 263.1176, 263.1176, 263.1176, 
    263.1176, 263.1176, 263.1176, 263.1176, 263.1176, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1172, 263.1172, 263.1172, 263.1172, 263.1172, 
    263.1172, 263.1173, 263.1174, 263.1173, 263.1174, 263.1174, 263.1174, 
    263.1174, 263.1174, 263.1175, 263.1174, 263.1176, 263.1175, 263.1176, 
    263.1176, 263.1176, 263.1176, 263.1177, 263.1177, 263.1177, 263.1178, 
    263.1172, 263.1172, 263.1172, 263.1173, 263.1173, 263.1174, 263.1175, 
    263.1174, 263.1175, 263.1175, 263.1174, 263.1175, 263.1173, 263.1173, 
    263.1173, 263.1172, 263.1174, 263.1173, 263.1175, 263.1175, 263.1176, 
    263.1176, 263.1177, 263.1178, 263.1179, 263.118, 263.1173, 263.1172, 
    263.1173, 263.1173, 263.1174, 263.1175, 263.1175, 263.1175, 263.1175, 
    263.1176, 263.1175, 263.1176, 263.1173, 263.1174, 263.1172, 263.1173, 
    263.1173, 263.1173, 263.1174, 263.1174, 263.1175, 263.1175, 263.1178, 
    263.1176, 263.118, 263.1179, 263.1172, 263.1173, 263.1174, 263.1173, 
    263.1175, 263.1175, 263.1175, 263.1176, 263.1176, 263.1176, 263.1176, 
    263.1176, 263.1175, 263.1175, 263.1174, 263.1174, 263.1174, 263.1174, 
    263.1174, 263.1175, 263.1175, 263.1175, 263.1176, 263.1175, 263.1178, 
    263.1176, 263.1173, 263.1174, 263.1174, 263.1173, 263.1175, 263.1175, 
    263.1176, 263.1176, 263.1176, 263.1176, 263.1176, 263.1176, 263.1175, 
    263.1175, 263.1174, 263.1173, 263.1174, 263.1174, 263.1175, 263.1176, 
    263.1176, 263.1176, 263.1175, 263.1175, 263.1175, 263.1176, 263.1174, 
    263.1176, 263.1174, 263.1174, 263.1175, 263.1175, 263.1176, 263.1176, 
    263.1176, 263.1175, 263.1175, 263.1174, 263.1174, 263.1174, 263.1174, 
    263.1174, 263.1174, 263.1175, 263.1176, 263.1176, 263.1176, 263.1177, 
    263.1177, 263.1178, 263.1177, 263.1179, 263.1176, 263.1177, 263.1175, 
    263.1175, 263.1175, 263.1176, 263.1176, 263.1176, 263.1175, 263.1174, 
    263.1174, 263.1174, 263.1174, 263.1174, 263.1174, 263.1174, 263.1175, 
    263.1175, 263.1176, 263.1176, 263.1178, 263.1179, 263.118, 263.118, 
    263.118, 263.118,
  263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.7253, 263.7362, 263.7341, 263.7429, 263.738, 263.7438, 263.7275, 
    263.7366, 263.7308, 263.7263, 263.7599, 263.7433, 263.7772, 263.7667, 
    263.7932, 263.7755, 263.7968, 263.7928, 263.805, 263.8015, 263.8171, 
    263.8066, 263.8252, 263.8146, 263.8163, 263.8063, 263.7467, 263.7578, 
    263.746, 263.7476, 263.7469, 263.7381, 263.7337, 263.7244, 263.7261, 
    263.7329, 263.7483, 263.7431, 263.7563, 263.756, 263.7706, 263.764, 
    263.7885, 263.7815, 263.8016, 263.7966, 263.8014, 263.7999, 263.8014, 
    263.794, 263.7972, 263.7906, 263.7652, 263.7726, 263.7503, 263.7368, 
    263.7279, 263.7215, 263.7224, 263.7241, 263.7329, 263.7412, 263.7476, 
    263.7518, 263.7559, 263.7684, 263.775, 263.7899, 263.7872, 263.7917, 
    263.7961, 263.8033, 263.8022, 263.8053, 263.7916, 263.8007, 263.7857, 
    263.7898, 263.757, 263.7445, 263.7391, 263.7345, 263.7231, 263.731, 
    263.7279, 263.7353, 263.7399, 263.7376, 263.7519, 263.7463, 263.7754, 
    263.7629, 263.7956, 263.7878, 263.7974, 263.7925, 263.801, 263.7934, 
    263.8065, 263.8094, 263.8074, 263.8149, 263.7929, 263.8014, 263.7375, 
    263.7379, 263.7397, 263.7319, 263.7315, 263.7244, 263.7307, 263.7334, 
    263.7402, 263.7442, 263.748, 263.7565, 263.7658, 263.7789, 263.7883, 
    263.7946, 263.7907, 263.7941, 263.7903, 263.7885, 263.8083, 263.7972, 
    263.8139, 263.813, 263.8054, 263.813, 263.7382, 263.736, 263.7285, 
    263.7344, 263.7236, 263.7296, 263.7331, 263.7464, 263.7494, 263.7521, 
    263.7575, 263.7643, 263.7763, 263.7868, 263.7963, 263.7956, 263.7959, 
    263.798, 263.7927, 263.7989, 263.7999, 263.7972, 263.8128, 263.8084, 
    263.8129, 263.81, 263.7367, 263.7404, 263.7384, 263.7421, 263.7395, 
    263.7511, 263.7546, 263.7708, 263.7642, 263.7747, 263.7653, 263.767, 
    263.7751, 263.7658, 263.7862, 263.7723, 263.7981, 263.7842, 263.799, 
    263.7963, 263.8007, 263.8047, 263.8096, 263.8188, 263.8167, 263.8243, 
    263.7458, 263.7505, 263.7502, 263.7551, 263.7588, 263.7667, 263.7793, 
    263.7745, 263.7833, 263.7851, 263.7718, 263.7799, 263.7537, 263.758, 
    263.7554, 263.7462, 263.7756, 263.7606, 263.7884, 263.7802, 263.8041, 
    263.7922, 263.8155, 263.8254, 263.8347, 263.8456, 263.7531, 263.7499, 
    263.7557, 263.7636, 263.7709, 263.7807, 263.7817, 263.7836, 263.7883, 
    263.7923, 263.7841, 263.7933, 263.7589, 263.7769, 263.7487, 263.7572, 
    263.7632, 263.7606, 263.774, 263.7772, 263.79, 263.7834, 263.8229, 
    263.8055, 263.8539, 263.8404, 263.7488, 263.7531, 263.7682, 263.761, 
    263.7814, 263.7864, 263.7905, 263.7957, 263.7963, 263.7993, 263.7943, 
    263.7992, 263.7808, 263.789, 263.7665, 263.7719, 263.7694, 263.7667, 
    263.7752, 263.7843, 263.7845, 263.7874, 263.7956, 263.7815, 263.8251, 
    263.7982, 263.7578, 263.7661, 263.7674, 263.7642, 263.7859, 263.778, 
    263.7993, 263.7935, 263.8029, 263.7983, 263.7976, 263.7916, 263.7878, 
    263.7784, 263.7707, 263.7646, 263.7661, 263.7727, 263.7848, 263.7963, 
    263.7938, 263.8022, 263.7799, 263.7893, 263.7856, 263.7951, 263.7744, 
    263.792, 263.77, 263.7719, 263.7778, 263.7899, 263.7926, 263.7954, 
    263.7937, 263.7851, 263.7838, 263.7777, 263.776, 263.7714, 263.7677, 
    263.7711, 263.7747, 263.7852, 263.7945, 263.8047, 263.8072, 263.819, 
    263.8094, 263.8253, 263.8117, 263.8352, 263.793, 263.8114, 263.7781, 
    263.7817, 263.7882, 263.803, 263.795, 263.8044, 263.7837, 263.7729, 
    263.7702, 263.765, 263.7703, 263.7699, 263.7749, 263.7733, 263.7855, 
    263.7789, 263.7976, 263.8044, 263.8235, 263.8352, 263.8471, 263.8524, 
    263.854, 263.8546 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  254.011, 254.0118, 254.0116, 254.0123, 254.0119, 254.0123, 254.0111, 
    254.0118, 254.0114, 254.011, 254.0135, 254.0123, 254.0148, 254.014, 
    254.016, 254.0147, 254.0163, 254.016, 254.0169, 254.0166, 254.0178, 
    254.017, 254.0184, 254.0176, 254.0177, 254.017, 254.0125, 254.0133, 
    254.0125, 254.0126, 254.0126, 254.0119, 254.0116, 254.0109, 254.011, 
    254.0115, 254.0127, 254.0123, 254.0133, 254.0132, 254.0143, 254.0138, 
    254.0157, 254.0151, 254.0166, 254.0163, 254.0166, 254.0165, 254.0166, 
    254.0161, 254.0163, 254.0158, 254.0139, 254.0145, 254.0128, 254.0118, 
    254.0112, 254.0107, 254.0108, 254.0109, 254.0115, 254.0121, 254.0126, 
    254.0129, 254.0132, 254.0141, 254.0146, 254.0157, 254.0156, 254.0159, 
    254.0162, 254.0168, 254.0167, 254.0169, 254.0159, 254.0166, 254.0154, 
    254.0157, 254.0133, 254.0124, 254.012, 254.0116, 254.0108, 254.0114, 
    254.0112, 254.0117, 254.0121, 254.0119, 254.0129, 254.0125, 254.0147, 
    254.0137, 254.0162, 254.0156, 254.0163, 254.016, 254.0166, 254.016, 
    254.017, 254.0172, 254.0171, 254.0176, 254.016, 254.0166, 254.0119, 
    254.0119, 254.012, 254.0115, 254.0114, 254.0109, 254.0114, 254.0116, 
    254.0121, 254.0124, 254.0126, 254.0133, 254.0139, 254.0149, 254.0156, 
    254.0161, 254.0158, 254.0161, 254.0158, 254.0157, 254.0171, 254.0163, 
    254.0175, 254.0175, 254.0169, 254.0175, 254.0119, 254.0118, 254.0112, 
    254.0116, 254.0108, 254.0113, 254.0115, 254.0125, 254.0128, 254.013, 
    254.0134, 254.0139, 254.0147, 254.0155, 254.0162, 254.0162, 254.0162, 
    254.0164, 254.016, 254.0164, 254.0165, 254.0163, 254.0175, 254.0171, 
    254.0175, 254.0173, 254.0118, 254.0121, 254.0119, 254.0122, 254.012, 
    254.0129, 254.0131, 254.0143, 254.0138, 254.0146, 254.0139, 254.014, 
    254.0146, 254.014, 254.0155, 254.0144, 254.0164, 254.0153, 254.0164, 
    254.0162, 254.0166, 254.0169, 254.0172, 254.0179, 254.0177, 254.0183, 
    254.0125, 254.0128, 254.0128, 254.0132, 254.0134, 254.014, 254.015, 
    254.0146, 254.0153, 254.0154, 254.0144, 254.015, 254.0131, 254.0134, 
    254.0132, 254.0125, 254.0147, 254.0136, 254.0156, 254.015, 254.0168, 
    254.0159, 254.0177, 254.0184, 254.0191, 254.0199, 254.013, 254.0128, 
    254.0132, 254.0138, 254.0143, 254.0151, 254.0152, 254.0153, 254.0156, 
    254.0159, 254.0153, 254.016, 254.0134, 254.0148, 254.0127, 254.0133, 
    254.0138, 254.0136, 254.0146, 254.0148, 254.0158, 254.0153, 254.0182, 
    254.0169, 254.0206, 254.0195, 254.0127, 254.013, 254.0141, 254.0136, 
    254.0151, 254.0155, 254.0158, 254.0162, 254.0162, 254.0165, 254.0161, 
    254.0164, 254.0151, 254.0157, 254.014, 254.0144, 254.0142, 254.014, 
    254.0147, 254.0153, 254.0154, 254.0156, 254.0161, 254.0151, 254.0183, 
    254.0163, 254.0134, 254.014, 254.0141, 254.0138, 254.0155, 254.0149, 
    254.0165, 254.016, 254.0167, 254.0164, 254.0163, 254.0159, 254.0156, 
    254.0149, 254.0143, 254.0139, 254.014, 254.0145, 254.0154, 254.0162, 
    254.016, 254.0167, 254.015, 254.0157, 254.0154, 254.0161, 254.0146, 
    254.0159, 254.0143, 254.0144, 254.0149, 254.0157, 254.016, 254.0162, 
    254.016, 254.0154, 254.0153, 254.0148, 254.0147, 254.0144, 254.0141, 
    254.0144, 254.0146, 254.0154, 254.0161, 254.0169, 254.0171, 254.0179, 
    254.0172, 254.0183, 254.0173, 254.0191, 254.016, 254.0173, 254.0149, 
    254.0152, 254.0156, 254.0167, 254.0161, 254.0168, 254.0153, 254.0145, 
    254.0143, 254.0139, 254.0143, 254.0143, 254.0146, 254.0145, 254.0154, 
    254.0149, 254.0163, 254.0168, 254.0183, 254.0191, 254.0201, 254.0204, 
    254.0206, 254.0206 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.1410976, 0.1411059, 0.1411043, 0.141111, 0.1411074, 0.1411116, 0.1410994, 
    0.1411062, 0.1411019, 0.1410985, 0.1411236, 0.1411113, 0.1411372, 
    0.1411292, 0.1411496, 0.1411358, 0.1411524, 0.1411493, 0.1411589, 
    0.1411562, 0.141168, 0.1411601, 0.1411744, 0.1411662, 0.1411674, 
    0.1411598, 0.1411139, 0.141122, 0.1411134, 0.1411146, 0.1411141, 
    0.1411074, 0.1411038, 0.1410971, 0.1410984, 0.1411034, 0.1411151, 
    0.1411112, 0.1411213, 0.1411211, 0.1411322, 0.1411272, 0.141146, 
    0.1411407, 0.1411563, 0.1411523, 0.1411561, 0.1411549, 0.1411561, 
    0.1411503, 0.1411528, 0.1411477, 0.1411281, 0.1411338, 0.1411167, 
    0.1411062, 0.1410996, 0.1410949, 0.1410955, 0.1410968, 0.1411034, 
    0.1411098, 0.1411147, 0.1411179, 0.141121, 0.1411302, 0.1411355, 
    0.141147, 0.1411451, 0.1411485, 0.1411519, 0.1411575, 0.1411566, 
    0.1411591, 0.1411485, 0.1411555, 0.141144, 0.1411471, 0.1411213, 
    0.1411123, 0.1411079, 0.1411046, 0.141096, 0.1411019, 0.1410996, 
    0.1411053, 0.1411088, 0.1411071, 0.1411179, 0.1411137, 0.1411358, 
    0.1411263, 0.1411515, 0.1411455, 0.141153, 0.1411492, 0.1411557, 
    0.1411499, 0.14116, 0.1411622, 0.1411607, 0.1411666, 0.1411495, 0.141156, 
    0.141107, 0.1411073, 0.1411086, 0.1411027, 0.1411023, 0.141097, 
    0.1411018, 0.1411038, 0.1411091, 0.1411121, 0.141115, 0.1411214, 
    0.1411285, 0.1411386, 0.1411459, 0.1411508, 0.1411478, 0.1411504, 
    0.1411475, 0.1411462, 0.1411613, 0.1411527, 0.1411657, 0.141165, 
    0.1411591, 0.1411651, 0.1411075, 0.1411059, 0.1411001, 0.1411046, 
    0.1410965, 0.1411009, 0.1411035, 0.1411137, 0.141116, 0.1411181, 
    0.1411222, 0.1411274, 0.1411366, 0.1411447, 0.1411522, 0.1411516, 
    0.1411518, 0.1411534, 0.1411494, 0.1411541, 0.1411548, 0.1411528, 
    0.1411649, 0.1411615, 0.141165, 0.1411628, 0.1411064, 0.1411092, 
    0.1411077, 0.1411105, 0.1411084, 0.1411172, 0.1411198, 0.1411323, 
    0.1411273, 0.1411354, 0.1411282, 0.1411294, 0.1411354, 0.1411286, 
    0.1411441, 0.1411334, 0.1411535, 0.1411425, 0.1411542, 0.1411521, 
    0.1411556, 0.1411586, 0.1411625, 0.1411695, 0.1411679, 0.1411738, 
    0.1411133, 0.1411168, 0.1411166, 0.1411204, 0.1411231, 0.1411293, 
    0.141139, 0.1411353, 0.1411421, 0.1411434, 0.1411332, 0.1411394, 
    0.1411193, 0.1411224, 0.1411206, 0.1411135, 0.141136, 0.1411244, 
    0.141146, 0.1411397, 0.1411581, 0.1411488, 0.141167, 0.1411744, 0.141182, 
    0.1411903, 0.1411189, 0.1411165, 0.1411209, 0.1411267, 0.1411325, 
    0.1411401, 0.1411409, 0.1411423, 0.141146, 0.1411491, 0.1411426, 
    0.1411498, 0.1411229, 0.1411371, 0.1411155, 0.1411218, 0.1411265, 
    0.1411245, 0.141135, 0.1411374, 0.1411472, 0.1411422, 0.1411725, 
    0.141159, 0.1411969, 0.1411862, 0.1411156, 0.1411189, 0.1411303, 
    0.1411249, 0.1411406, 0.1411445, 0.1411477, 0.1411516, 0.1411521, 
    0.1411545, 0.1411506, 0.1411543, 0.1411401, 0.1411465, 0.1411291, 
    0.1411333, 0.1411314, 0.1411293, 0.1411359, 0.1411427, 0.141143, 
    0.1411452, 0.1411509, 0.1411407, 0.1411739, 0.141153, 0.1411225, 
    0.1411286, 0.1411297, 0.1411273, 0.1411441, 0.141138, 0.1411544, 0.14115, 
    0.1411573, 0.1411537, 0.1411531, 0.1411485, 0.1411456, 0.1411382, 
    0.1411323, 0.1411277, 0.1411288, 0.1411338, 0.1411431, 0.1411521, 
    0.1411501, 0.1411567, 0.1411395, 0.1411466, 0.1411438, 0.1411512, 
    0.1411352, 0.1411482, 0.1411318, 0.1411333, 0.1411379, 0.141147, 
    0.1411493, 0.1411514, 0.1411501, 0.1411434, 0.1411424, 0.1411378, 
    0.1411364, 0.141133, 0.14113, 0.1411327, 0.1411354, 0.1411435, 0.1411507, 
    0.1411586, 0.1411606, 0.1411694, 0.141162, 0.1411739, 0.1411634, 
    0.1411819, 0.1411493, 0.1411634, 0.1411381, 0.1411409, 0.1411457, 
    0.1411571, 0.1411512, 0.1411582, 0.1411424, 0.1411339, 0.141132, 
    0.1411279, 0.1411321, 0.1411317, 0.1411357, 0.1411344, 0.1411438, 
    0.1411387, 0.1411531, 0.1411582, 0.1411731, 0.1411822, 0.1411917, 
    0.1411958, 0.1411971, 0.1411976,
  0.147692, 0.1477012, 0.1476994, 0.1477067, 0.1477027, 0.1477075, 0.147694, 
    0.1477015, 0.1476967, 0.147693, 0.1477206, 0.1477071, 0.1477356, 
    0.1477268, 0.1477492, 0.1477341, 0.1477523, 0.147749, 0.1477595, 
    0.1477565, 0.1477696, 0.1477609, 0.1477767, 0.1477676, 0.1477689, 
    0.1477606, 0.14771, 0.1477189, 0.1477094, 0.1477107, 0.1477101, 
    0.1477028, 0.1476989, 0.1476915, 0.1476928, 0.1476984, 0.1477113, 
    0.147707, 0.1477181, 0.1477178, 0.1477301, 0.1477246, 0.1477453, 
    0.1477395, 0.1477566, 0.1477523, 0.1477564, 0.1477551, 0.1477564, 
    0.14775, 0.1477527, 0.1477472, 0.1477256, 0.1477319, 0.147713, 0.1477015, 
    0.1476943, 0.147689, 0.1476898, 0.1476911, 0.1476984, 0.1477055, 
    0.1477108, 0.1477143, 0.1477178, 0.147728, 0.1477337, 0.1477464, 
    0.1477443, 0.147748, 0.1477518, 0.147758, 0.147757, 0.1477597, 0.1477481, 
    0.1477557, 0.147743, 0.1477465, 0.1477181, 0.1477082, 0.1477034, 
    0.1476997, 0.1476903, 0.1476968, 0.1476942, 0.1477005, 0.1477043, 
    0.1477025, 0.1477144, 0.1477097, 0.1477341, 0.1477236, 0.1477514, 
    0.1477447, 0.147753, 0.1477488, 0.147756, 0.1477495, 0.1477608, 
    0.1477631, 0.1477615, 0.147768, 0.1477492, 0.1477563, 0.1477024, 
    0.1477027, 0.1477042, 0.1476976, 0.1476972, 0.1476914, 0.1476966, 
    0.1476988, 0.1477046, 0.1477079, 0.1477111, 0.1477182, 0.147726, 
    0.1477371, 0.1477452, 0.1477506, 0.1477473, 0.1477502, 0.1477469, 
    0.1477454, 0.1477622, 0.1477527, 0.1477671, 0.1477663, 0.1477598, 
    0.1477664, 0.1477029, 0.1477011, 0.1476948, 0.1476997, 0.1476908, 
    0.1476957, 0.1476985, 0.1477097, 0.1477123, 0.1477145, 0.1477191, 
    0.1477248, 0.1477349, 0.1477438, 0.1477521, 0.1477515, 0.1477517, 
    0.1477535, 0.147749, 0.1477542, 0.147755, 0.1477528, 0.1477662, 
    0.1477624, 0.1477663, 0.1477638, 0.1477017, 0.1477047, 0.1477031, 
    0.1477062, 0.1477039, 0.1477136, 0.1477164, 0.1477302, 0.1477247, 
    0.1477336, 0.1477256, 0.147727, 0.1477336, 0.1477261, 0.1477432, 
    0.1477314, 0.1477535, 0.1477414, 0.1477543, 0.147752, 0.1477558, 
    0.1477591, 0.1477634, 0.1477712, 0.1477694, 0.147776, 0.1477093, 
    0.1477132, 0.1477129, 0.1477171, 0.1477201, 0.1477268, 0.1477375, 
    0.1477335, 0.147741, 0.1477424, 0.1477312, 0.147738, 0.1477159, 
    0.1477193, 0.1477173, 0.1477095, 0.1477343, 0.1477215, 0.1477453, 
    0.1477384, 0.1477586, 0.1477484, 0.1477684, 0.1477767, 0.147785, 
    0.1477942, 0.1477154, 0.1477128, 0.1477176, 0.1477241, 0.1477305, 
    0.1477388, 0.1477397, 0.1477412, 0.1477453, 0.1477486, 0.1477416, 
    0.1477495, 0.1477199, 0.1477355, 0.1477117, 0.1477187, 0.1477238, 
    0.1477216, 0.1477331, 0.1477358, 0.1477466, 0.1477411, 0.1477745, 
    0.1477597, 0.1478016, 0.1477897, 0.1477118, 0.1477154, 0.147728, 
    0.147722, 0.1477394, 0.1477436, 0.1477471, 0.1477515, 0.147752, 
    0.1477546, 0.1477504, 0.1477545, 0.1477388, 0.1477458, 0.1477267, 
    0.1477313, 0.1477292, 0.1477268, 0.1477341, 0.1477416, 0.147742, 
    0.1477444, 0.1477508, 0.1477394, 0.1477761, 0.1477531, 0.1477194, 
    0.1477262, 0.1477274, 0.1477247, 0.1477432, 0.1477364, 0.1477546, 
    0.1477497, 0.1477577, 0.1477537, 0.1477531, 0.147748, 0.1477448, 
    0.1477367, 0.1477302, 0.1477251, 0.1477263, 0.1477319, 0.1477421, 
    0.147752, 0.1477498, 0.1477571, 0.1477381, 0.147746, 0.1477429, 0.147751, 
    0.1477334, 0.1477478, 0.1477297, 0.1477313, 0.1477363, 0.1477464, 
    0.1477489, 0.1477512, 0.1477498, 0.1477424, 0.1477413, 0.1477362, 
    0.1477347, 0.1477309, 0.1477277, 0.1477306, 0.1477336, 0.1477425, 
    0.1477504, 0.1477592, 0.1477614, 0.1477711, 0.1477629, 0.1477762, 
    0.1477645, 0.147785, 0.1477489, 0.1477646, 0.1477366, 0.1477396, 
    0.147745, 0.1477576, 0.147751, 0.1477588, 0.1477413, 0.147732, 0.1477298, 
    0.1477254, 0.1477299, 0.1477296, 0.1477339, 0.1477325, 0.1477428, 
    0.1477373, 0.1477531, 0.1477588, 0.1477752, 0.1477853, 0.1477958, 
    0.1478003, 0.1478017, 0.1478023,
  0.1573315, 0.157342, 0.15734, 0.1573484, 0.1573438, 0.1573493, 0.1573337, 
    0.1573424, 0.1573369, 0.1573326, 0.1573646, 0.1573488, 0.1573818, 
    0.1573715, 0.1573975, 0.1573801, 0.1574011, 0.1573972, 0.1574093, 
    0.1574058, 0.1574211, 0.1574109, 0.1574292, 0.1574187, 0.1574203, 
    0.1574105, 0.1573522, 0.1573626, 0.1573515, 0.157353, 0.1573524, 
    0.1573439, 0.1573395, 0.1573308, 0.1573324, 0.1573389, 0.1573537, 
    0.1573487, 0.1573615, 0.1573612, 0.1573754, 0.157369, 0.157393, 
    0.1573862, 0.157406, 0.157401, 0.1574057, 0.1574043, 0.1574057, 
    0.1573984, 0.1574015, 0.1573951, 0.1573701, 0.1573774, 0.1573557, 
    0.1573424, 0.1573341, 0.157328, 0.1573289, 0.1573305, 0.1573389, 
    0.1573469, 0.1573531, 0.1573571, 0.1573612, 0.157373, 0.1573796, 
    0.1573942, 0.1573918, 0.1573961, 0.1574005, 0.1574076, 0.1574065, 
    0.1574096, 0.1573961, 0.157405, 0.1573903, 0.1573943, 0.1573617, 
    0.1573501, 0.1573447, 0.1573404, 0.1573295, 0.157337, 0.157334, 
    0.1573412, 0.1573457, 0.1573435, 0.1573572, 0.1573519, 0.15738, 
    0.1573679, 0.1574, 0.1573923, 0.1574018, 0.157397, 0.1574052, 0.1573978, 
    0.1574108, 0.1574136, 0.1574116, 0.1574192, 0.1573974, 0.1574057, 
    0.1573434, 0.1573437, 0.1573455, 0.1573379, 0.1573375, 0.1573308, 
    0.1573368, 0.1573393, 0.157346, 0.1573498, 0.1573535, 0.1573616, 
    0.1573707, 0.1573835, 0.1573928, 0.157399, 0.1573952, 0.1573986, 
    0.1573948, 0.1573931, 0.1574125, 0.1574015, 0.1574181, 0.1574172, 
    0.1574096, 0.1574173, 0.157344, 0.157342, 0.1573347, 0.1573404, 0.15733, 
    0.1573357, 0.157339, 0.1573519, 0.1573548, 0.1573574, 0.1573626, 
    0.1573693, 0.157381, 0.1573913, 0.1574007, 0.1574001, 0.1574003, 
    0.1574024, 0.1573972, 0.1574032, 0.1574042, 0.1574016, 0.1574171, 
    0.1574126, 0.1574172, 0.1574143, 0.1573426, 0.1573461, 0.1573442, 
    0.1573478, 0.1573452, 0.1573563, 0.1573597, 0.1573755, 0.1573691, 
    0.1573794, 0.1573702, 0.1573718, 0.1573795, 0.1573707, 0.1573906, 
    0.1573769, 0.1574024, 0.1573885, 0.1574033, 0.1574007, 0.1574051, 
    0.1574089, 0.1574139, 0.1574229, 0.1574208, 0.1574284, 0.1573514, 
    0.1573559, 0.1573556, 0.1573603, 0.1573638, 0.1573716, 0.1573839, 
    0.1573793, 0.1573879, 0.1573896, 0.1573766, 0.1573845, 0.1573589, 
    0.157363, 0.1573606, 0.1573517, 0.1573803, 0.1573655, 0.1573929, 
    0.1573849, 0.1574083, 0.1573966, 0.1574197, 0.1574293, 0.1574389, 
    0.1574496, 0.1573584, 0.1573554, 0.1573609, 0.1573685, 0.1573758, 
    0.1573854, 0.1573864, 0.1573882, 0.1573929, 0.1573968, 0.1573886, 
    0.1573978, 0.1573637, 0.1573816, 0.1573541, 0.1573622, 0.1573681, 
    0.1573656, 0.1573788, 0.1573819, 0.1573945, 0.157388, 0.1574268, 
    0.1574096, 0.1574581, 0.1574444, 0.1573543, 0.1573585, 0.157373, 
    0.1573661, 0.157386, 0.1573909, 0.157395, 0.1574001, 0.1574007, 
    0.1574037, 0.1573987, 0.1574035, 0.1573854, 0.1573935, 0.1573714, 
    0.1573767, 0.1573743, 0.1573716, 0.15738, 0.1573887, 0.1573891, 
    0.1573919, 0.1573994, 0.1573862, 0.1574287, 0.1574021, 0.157363, 
    0.1573709, 0.1573722, 0.1573691, 0.1573904, 0.1573827, 0.1574036, 
    0.157398, 0.1574073, 0.1574026, 0.157402, 0.1573961, 0.1573924, 0.157383, 
    0.1573755, 0.1573696, 0.157371, 0.1573775, 0.1573893, 0.1574007, 
    0.1573981, 0.1574066, 0.1573846, 0.1573937, 0.1573901, 0.1573995, 
    0.1573792, 0.157396, 0.1573748, 0.1573767, 0.1573825, 0.1573942, 
    0.1573971, 0.1573998, 0.1573981, 0.1573896, 0.1573883, 0.1573824, 
    0.1573807, 0.1573763, 0.1573726, 0.157376, 0.1573795, 0.1573897, 
    0.1573989, 0.1574089, 0.1574115, 0.1574229, 0.1574134, 0.1574288, 
    0.1574153, 0.1574389, 0.1573972, 0.1574153, 0.1573829, 0.1573864, 
    0.1573926, 0.1574072, 0.1573995, 0.1574086, 0.1573883, 0.1573776, 
    0.157375, 0.1573699, 0.1573752, 0.1573747, 0.1573797, 0.1573781, 0.15739, 
    0.1573837, 0.1574019, 0.1574085, 0.1574276, 0.1574392, 0.1574513, 
    0.1574566, 0.1574582, 0.1574589,
  0.1706156, 0.170627, 0.1706248, 0.170634, 0.170629, 0.170635, 0.170618, 
    0.1706274, 0.1706214, 0.1706167, 0.1706518, 0.1706345, 0.1706704, 
    0.1706592, 0.1706876, 0.1706686, 0.1706914, 0.1706871, 0.1707004, 
    0.1706966, 0.1707133, 0.1707021, 0.1707222, 0.1707107, 0.1707125, 
    0.1707017, 0.1706381, 0.1706496, 0.1706373, 0.170639, 0.1706383, 
    0.170629, 0.1706243, 0.1706148, 0.1706166, 0.1706236, 0.1706397, 
    0.1706343, 0.1706482, 0.1706479, 0.1706633, 0.1706564, 0.1706825, 
    0.1706751, 0.1706967, 0.1706913, 0.1706965, 0.1706949, 0.1706965, 
    0.1706885, 0.1706919, 0.1706849, 0.1706576, 0.1706656, 0.1706419, 
    0.1706276, 0.1706184, 0.1706118, 0.1706127, 0.1706145, 0.1706236, 
    0.1706324, 0.170639, 0.1706434, 0.1706479, 0.1706609, 0.1706681, 
    0.170684, 0.1706812, 0.170686, 0.1706907, 0.1706985, 0.1706973, 
    0.1707007, 0.170686, 0.1706957, 0.1706796, 0.170684, 0.1706486, 
    0.1706358, 0.17063, 0.1706253, 0.1706134, 0.1706215, 0.1706183, 
    0.1706261, 0.170631, 0.1706286, 0.1706436, 0.1706377, 0.1706685, 
    0.1706552, 0.1706902, 0.1706818, 0.1706922, 0.1706869, 0.170696, 
    0.1706878, 0.170702, 0.1707051, 0.170703, 0.1707111, 0.1706874, 
    0.1706964, 0.1706285, 0.1706289, 0.1706307, 0.1706226, 0.1706221, 
    0.1706147, 0.1706213, 0.1706241, 0.1706313, 0.1706355, 0.1706395, 
    0.1706484, 0.1706582, 0.1706722, 0.1706823, 0.1706891, 0.170685, 
    0.1706886, 0.1706845, 0.1706826, 0.1707039, 0.1706919, 0.17071, 0.170709, 
    0.1707008, 0.1707091, 0.1706292, 0.1706269, 0.170619, 0.1706252, 
    0.1706139, 0.1706202, 0.1706237, 0.1706377, 0.1706409, 0.1706438, 
    0.1706495, 0.1706567, 0.1706695, 0.1706807, 0.170691, 0.1706903, 
    0.1706905, 0.1706928, 0.1706871, 0.1706937, 0.1706948, 0.170692, 
    0.1707089, 0.170704, 0.170709, 0.1707058, 0.1706277, 0.1706315, 
    0.1706294, 0.1706333, 0.1706305, 0.1706426, 0.1706463, 0.1706635, 
    0.1706566, 0.1706678, 0.1706577, 0.1706595, 0.170668, 0.1706583, 0.17068, 
    0.1706651, 0.1706929, 0.1706778, 0.1706938, 0.170691, 0.1706958, 0.1707, 
    0.1707054, 0.1707152, 0.170713, 0.1707213, 0.1706372, 0.1706421, 
    0.1706418, 0.170647, 0.1706508, 0.1706592, 0.1706727, 0.1706677, 
    0.170677, 0.1706789, 0.1706647, 0.1706733, 0.1706455, 0.1706499, 
    0.1706473, 0.1706375, 0.1706687, 0.1706526, 0.1706825, 0.1706737, 
    0.1706994, 0.1706865, 0.1707117, 0.1707223, 0.1707327, 0.1707445, 
    0.1706449, 0.1706415, 0.1706476, 0.1706559, 0.1706638, 0.1706742, 
    0.1706754, 0.1706773, 0.1706824, 0.1706867, 0.1706779, 0.1706878, 
    0.1706507, 0.1706702, 0.1706402, 0.1706491, 0.1706554, 0.1706527, 
    0.1706671, 0.1706705, 0.1706842, 0.1706772, 0.1707196, 0.1707008, 
    0.1707538, 0.1707388, 0.1706403, 0.1706449, 0.1706607, 0.1706532, 
    0.170675, 0.1706803, 0.1706848, 0.1706903, 0.170691, 0.1706943, 
    0.1706889, 0.1706941, 0.1706743, 0.1706831, 0.170659, 0.1706648, 
    0.1706622, 0.1706592, 0.1706683, 0.170678, 0.1706783, 0.1706814, 
    0.1706898, 0.1706751, 0.1707218, 0.1706927, 0.1706499, 0.1706585, 
    0.1706599, 0.1706565, 0.1706798, 0.1706713, 0.1706942, 0.170688, 
    0.1706982, 0.1706931, 0.1706924, 0.1706859, 0.1706819, 0.1706717, 
    0.1706635, 0.1706571, 0.1706586, 0.1706656, 0.1706786, 0.170691, 
    0.1706882, 0.1706974, 0.1706734, 0.1706834, 0.1706795, 0.1706897, 
    0.1706675, 0.170686, 0.1706627, 0.1706648, 0.1706712, 0.170684, 0.170687, 
    0.17069, 0.1706882, 0.1706789, 0.1706775, 0.1706711, 0.1706692, 
    0.1706644, 0.1706603, 0.170664, 0.1706678, 0.170679, 0.170689, 0.1707, 
    0.1707028, 0.1707153, 0.1707049, 0.170722, 0.1707072, 0.170733, 
    0.1706873, 0.170707, 0.1706715, 0.1706754, 0.1706822, 0.1706981, 
    0.1706896, 0.1706996, 0.1706774, 0.1706658, 0.170663, 0.1706574, 
    0.1706631, 0.1706626, 0.1706681, 0.1706663, 0.1706794, 0.1706724, 
    0.1706923, 0.1706996, 0.1707204, 0.1707331, 0.1707464, 0.1707522, 
    0.1707539, 0.1707547,
  0.1854066, 0.1854161, 0.1854143, 0.1854219, 0.1854177, 0.1854227, 
    0.1854085, 0.1854164, 0.1854114, 0.1854075, 0.1854368, 0.1854223, 
    0.1854522, 0.1854428, 0.1854665, 0.1854507, 0.1854697, 0.1854661, 
    0.1854772, 0.185474, 0.185488, 0.1854786, 0.1854954, 0.1854858, 
    0.1854873, 0.1854783, 0.1854252, 0.1854349, 0.1854247, 0.185426, 
    0.1854254, 0.1854178, 0.1854139, 0.1854059, 0.1854074, 0.1854132, 
    0.1854267, 0.1854221, 0.1854337, 0.1854334, 0.1854463, 0.1854405, 
    0.1854623, 0.1854561, 0.1854741, 0.1854696, 0.1854739, 0.1854726, 
    0.1854739, 0.1854672, 0.1854701, 0.1854642, 0.1854416, 0.1854482, 
    0.1854284, 0.1854166, 0.1854089, 0.1854034, 0.1854042, 0.1854056, 
    0.1854133, 0.1854205, 0.185426, 0.1854297, 0.1854334, 0.1854443, 
    0.1854503, 0.1854635, 0.1854612, 0.1854652, 0.1854691, 0.1854756, 
    0.1854746, 0.1854774, 0.1854651, 0.1854733, 0.1854598, 0.1854635, 
    0.1854341, 0.1854234, 0.1854186, 0.1854146, 0.1854048, 0.1854115, 
    0.1854089, 0.1854153, 0.1854194, 0.1854174, 0.1854298, 0.185425, 
    0.1854506, 0.1854395, 0.1854686, 0.1854617, 0.1854703, 0.1854659, 
    0.1854735, 0.1854667, 0.1854785, 0.1854811, 0.1854793, 0.1854862, 
    0.1854663, 0.1854739, 0.1854173, 0.1854176, 0.1854191, 0.1854124, 
    0.185412, 0.1854059, 0.1854113, 0.1854136, 0.1854196, 0.1854231, 
    0.1854265, 0.1854338, 0.1854421, 0.1854537, 0.1854621, 0.1854678, 
    0.1854643, 0.1854674, 0.185464, 0.1854624, 0.1854801, 0.1854701, 
    0.1854852, 0.1854843, 0.1854775, 0.1854844, 0.1854178, 0.185416, 
    0.1854094, 0.1854145, 0.1854052, 0.1854104, 0.1854134, 0.185425, 
    0.1854276, 0.18543, 0.1854347, 0.1854408, 0.1854514, 0.1854608, 
    0.1854694, 0.1854687, 0.1854689, 0.1854708, 0.1854661, 0.1854716, 
    0.1854725, 0.1854701, 0.1854842, 0.1854802, 0.1854843, 0.1854817, 
    0.1854166, 0.1854198, 0.185418, 0.1854213, 0.185419, 0.1854291, 
    0.1854322, 0.1854465, 0.1854407, 0.18545, 0.1854416, 0.1854431, 
    0.1854502, 0.1854421, 0.1854602, 0.1854478, 0.1854709, 0.1854584, 
    0.1854717, 0.1854693, 0.1854733, 0.1854768, 0.1854813, 0.1854896, 
    0.1854877, 0.1854946, 0.1854245, 0.1854286, 0.1854283, 0.1854326, 
    0.1854358, 0.1854429, 0.1854541, 0.1854499, 0.1854577, 0.1854592, 
    0.1854474, 0.1854546, 0.1854314, 0.1854351, 0.1854329, 0.1854248, 
    0.1854508, 0.1854374, 0.1854623, 0.1854549, 0.1854763, 0.1854656, 
    0.1854866, 0.1854955, 0.1855042, 0.1855141, 0.1854309, 0.1854281, 
    0.1854332, 0.1854401, 0.1854467, 0.1854554, 0.1854563, 0.1854579, 
    0.1854622, 0.1854658, 0.1854584, 0.1854666, 0.1854359, 0.185452, 
    0.185427, 0.1854344, 0.1854397, 0.1854375, 0.1854494, 0.1854522, 
    0.1854637, 0.1854578, 0.1854933, 0.1854775, 0.1855218, 0.1855093, 
    0.1854271, 0.1854309, 0.1854441, 0.1854379, 0.185456, 0.1854605, 
    0.1854641, 0.1854688, 0.1854693, 0.1854721, 0.1854675, 0.1854719, 
    0.1854554, 0.1854628, 0.1854427, 0.1854475, 0.1854453, 0.1854428, 
    0.1854504, 0.1854585, 0.1854587, 0.1854613, 0.1854685, 0.1854561, 
    0.1854952, 0.1854709, 0.1854351, 0.1854423, 0.1854434, 0.1854406, 
    0.18546, 0.185453, 0.185472, 0.1854669, 0.1854753, 0.1854711, 0.1854705, 
    0.1854651, 0.1854617, 0.1854533, 0.1854464, 0.185441, 0.1854423, 
    0.1854482, 0.185459, 0.1854693, 0.185467, 0.1854747, 0.1854547, 0.185463, 
    0.1854598, 0.1854682, 0.1854498, 0.1854653, 0.1854458, 0.1854475, 
    0.1854528, 0.1854635, 0.185466, 0.1854685, 0.185467, 0.1854593, 
    0.1854581, 0.1854527, 0.1854512, 0.1854471, 0.1854437, 0.1854468, 
    0.1854501, 0.1854593, 0.1854677, 0.1854769, 0.1854791, 0.1854897, 
    0.185481, 0.1854953, 0.185483, 0.1855045, 0.1854663, 0.1854828, 
    0.1854531, 0.1854563, 0.185462, 0.1854753, 0.1854682, 0.1854766, 
    0.185458, 0.1854484, 0.185446, 0.1854414, 0.1854461, 0.1854457, 
    0.1854502, 0.1854488, 0.1854596, 0.1854538, 0.1854704, 0.1854765, 
    0.1854939, 0.1855046, 0.1855156, 0.1855204, 0.1855219, 0.1855225,
  0.1954522, 0.1954562, 0.1954554, 0.1954586, 0.1954568, 0.1954589, 0.195453, 
    0.1954563, 0.1954542, 0.1954525, 0.1954649, 0.1954588, 0.1954714, 
    0.1954675, 0.1954775, 0.1954708, 0.1954789, 0.1954773, 0.195482, 
    0.1954807, 0.1954866, 0.1954826, 0.1954898, 0.1954857, 0.1954863, 
    0.1954825, 0.19546, 0.1954641, 0.1954598, 0.1954604, 0.1954601, 
    0.1954569, 0.1954552, 0.1954519, 0.1954525, 0.195455, 0.1954606, 
    0.1954587, 0.1954636, 0.1954635, 0.1954689, 0.1954665, 0.1954757, 
    0.1954731, 0.1954807, 0.1954788, 0.1954806, 0.1954801, 0.1954806, 
    0.1954778, 0.195479, 0.1954765, 0.1954669, 0.1954697, 0.1954614, 
    0.1954564, 0.1954531, 0.1954508, 0.1954511, 0.1954518, 0.195455, 
    0.195458, 0.1954604, 0.1954619, 0.1954635, 0.1954681, 0.1954706, 
    0.1954762, 0.1954752, 0.1954769, 0.1954786, 0.1954814, 0.1954809, 
    0.1954821, 0.1954769, 0.1954804, 0.1954747, 0.1954762, 0.1954638, 
    0.1954592, 0.1954572, 0.1954555, 0.1954514, 0.1954542, 0.1954531, 
    0.1954558, 0.1954575, 0.1954567, 0.195462, 0.1954599, 0.1954708, 
    0.1954661, 0.1954784, 0.1954754, 0.1954791, 0.1954772, 0.1954805, 
    0.1954776, 0.1954826, 0.1954837, 0.1954829, 0.1954858, 0.1954774, 
    0.1954806, 0.1954567, 0.1954568, 0.1954574, 0.1954546, 0.1954544, 
    0.1954518, 0.1954542, 0.1954551, 0.1954577, 0.1954591, 0.1954605, 
    0.1954637, 0.1954672, 0.1954721, 0.1954756, 0.195478, 0.1954766, 
    0.1954779, 0.1954764, 0.1954757, 0.1954833, 0.195479, 0.1954854, 
    0.1954851, 0.1954822, 0.1954851, 0.1954569, 0.1954561, 0.1954533, 
    0.1954555, 0.1954516, 0.1954537, 0.195455, 0.1954599, 0.195461, 0.195462, 
    0.195464, 0.1954666, 0.1954711, 0.1954751, 0.1954787, 0.1954784, 
    0.1954785, 0.1954793, 0.1954773, 0.1954797, 0.19548, 0.195479, 0.195485, 
    0.1954833, 0.195485, 0.1954839, 0.1954564, 0.1954577, 0.195457, 
    0.1954583, 0.1954574, 0.1954617, 0.195463, 0.195469, 0.1954665, 
    0.1954705, 0.195467, 0.1954676, 0.1954706, 0.1954671, 0.1954748, 
    0.1954696, 0.1954794, 0.1954741, 0.1954797, 0.1954787, 0.1954804, 
    0.1954819, 0.1954838, 0.1954873, 0.1954865, 0.1954894, 0.1954597, 
    0.1954615, 0.1954613, 0.1954632, 0.1954645, 0.1954675, 0.1954722, 
    0.1954705, 0.1954737, 0.1954744, 0.1954694, 0.1954725, 0.1954626, 
    0.1954642, 0.1954633, 0.1954599, 0.1954708, 0.1954652, 0.1954757, 
    0.1954726, 0.1954816, 0.1954771, 0.195486, 0.1954898, 0.1954935, 
    0.1954977, 0.1954624, 0.1954612, 0.1954634, 0.1954663, 0.1954691, 
    0.1954728, 0.1954732, 0.1954738, 0.1954757, 0.1954772, 0.1954741, 
    0.1954775, 0.1954646, 0.1954713, 0.1954608, 0.1954639, 0.1954662, 
    0.1954652, 0.1954702, 0.1954714, 0.1954763, 0.1954738, 0.1954889, 
    0.1954822, 0.195501, 0.1954957, 0.1954608, 0.1954624, 0.195468, 
    0.1954654, 0.195473, 0.1954749, 0.1954765, 0.1954785, 0.1954787, 
    0.1954799, 0.1954779, 0.1954798, 0.1954728, 0.1954759, 0.1954674, 
    0.1954695, 0.1954685, 0.1954675, 0.1954707, 0.1954741, 0.1954742, 
    0.1954753, 0.1954784, 0.1954731, 0.1954897, 0.1954794, 0.1954642, 
    0.1954673, 0.1954677, 0.1954665, 0.1954747, 0.1954717, 0.1954798, 
    0.1954776, 0.1954812, 0.1954794, 0.1954792, 0.1954769, 0.1954755, 
    0.1954719, 0.195469, 0.1954667, 0.1954672, 0.1954698, 0.1954743, 
    0.1954787, 0.1954777, 0.1954809, 0.1954725, 0.195476, 0.1954746, 
    0.1954782, 0.1954704, 0.195477, 0.1954687, 0.1954694, 0.1954717, 
    0.1954762, 0.1954773, 0.1954783, 0.1954777, 0.1954744, 0.1954739, 
    0.1954716, 0.195471, 0.1954693, 0.1954678, 0.1954692, 0.1954705, 
    0.1954744, 0.195478, 0.1954819, 0.1954829, 0.1954874, 0.1954837, 
    0.1954898, 0.1954845, 0.1954936, 0.1954774, 0.1954844, 0.1954718, 
    0.1954732, 0.1954756, 0.1954812, 0.1954782, 0.1954818, 0.1954739, 
    0.1954698, 0.1954688, 0.1954668, 0.1954688, 0.1954687, 0.1954706, 
    0.19547, 0.1954746, 0.1954721, 0.1954792, 0.1954817, 0.1954891, 
    0.1954937, 0.1954983, 0.1955004, 0.195501, 0.1955013,
  0.1982578, 0.1982584, 0.1982583, 0.1982588, 0.1982585, 0.1982588, 
    0.1982579, 0.1982584, 0.1982581, 0.1982579, 0.1982597, 0.1982588, 
    0.1982607, 0.1982601, 0.1982616, 0.1982606, 0.1982618, 0.1982616, 
    0.1982623, 0.1982621, 0.198263, 0.1982624, 0.1982635, 0.1982629, 
    0.198263, 0.1982624, 0.198259, 0.1982596, 0.198259, 0.198259, 0.198259, 
    0.1982585, 0.1982583, 0.1982578, 0.1982579, 0.1982582, 0.1982591, 
    0.1982588, 0.1982595, 0.1982595, 0.1982603, 0.19826, 0.1982614, 0.198261, 
    0.1982621, 0.1982618, 0.1982621, 0.198262, 0.1982621, 0.1982617, 
    0.1982619, 0.1982615, 0.19826, 0.1982605, 0.1982592, 0.1982584, 0.198258, 
    0.1982576, 0.1982577, 0.1982577, 0.1982582, 0.1982587, 0.198259, 
    0.1982593, 0.1982595, 0.1982602, 0.1982606, 0.1982614, 0.1982613, 
    0.1982616, 0.1982618, 0.1982622, 0.1982622, 0.1982623, 0.1982615, 
    0.1982621, 0.1982612, 0.1982614, 0.1982596, 0.1982589, 0.1982586, 
    0.1982583, 0.1982577, 0.1982581, 0.198258, 0.1982584, 0.1982586, 
    0.1982585, 0.1982593, 0.198259, 0.1982606, 0.1982599, 0.1982618, 
    0.1982613, 0.1982619, 0.1982616, 0.1982621, 0.1982616, 0.1982624, 
    0.1982626, 0.1982625, 0.1982629, 0.1982616, 0.1982621, 0.1982585, 
    0.1982585, 0.1982586, 0.1982582, 0.1982581, 0.1982578, 0.1982581, 
    0.1982583, 0.1982586, 0.1982589, 0.1982591, 0.1982595, 0.1982601, 
    0.1982608, 0.1982614, 0.1982617, 0.1982615, 0.1982617, 0.1982615, 
    0.1982614, 0.1982625, 0.1982619, 0.1982628, 0.1982628, 0.1982623, 
    0.1982628, 0.1982585, 0.1982584, 0.198258, 0.1982583, 0.1982577, 
    0.1982581, 0.1982582, 0.198259, 0.1982591, 0.1982593, 0.1982596, 0.19826, 
    0.1982607, 0.1982613, 0.1982618, 0.1982618, 0.1982618, 0.1982619, 
    0.1982616, 0.198262, 0.198262, 0.1982619, 0.1982628, 0.1982625, 
    0.1982628, 0.1982626, 0.1982584, 0.1982586, 0.1982585, 0.1982587, 
    0.1982586, 0.1982592, 0.1982594, 0.1982604, 0.19826, 0.1982606, 0.19826, 
    0.1982601, 0.1982606, 0.1982601, 0.1982612, 0.1982604, 0.1982619, 
    0.1982611, 0.198262, 0.1982618, 0.1982621, 0.1982623, 0.1982626, 
    0.1982631, 0.198263, 0.1982635, 0.198259, 0.1982592, 0.1982592, 
    0.1982595, 0.1982597, 0.1982601, 0.1982608, 0.1982606, 0.1982611, 
    0.1982612, 0.1982604, 0.1982609, 0.1982594, 0.1982596, 0.1982595, 
    0.198259, 0.1982606, 0.1982598, 0.1982614, 0.1982609, 0.1982623, 
    0.1982616, 0.1982629, 0.1982635, 0.1982641, 0.1982647, 0.1982594, 
    0.1982592, 0.1982595, 0.1982599, 0.1982604, 0.1982609, 0.198261, 
    0.1982611, 0.1982614, 0.1982616, 0.1982611, 0.1982616, 0.1982597, 
    0.1982607, 0.1982591, 0.1982596, 0.1982599, 0.1982598, 0.1982605, 
    0.1982607, 0.1982615, 0.1982611, 0.1982634, 0.1982623, 0.1982652, 
    0.1982644, 0.1982591, 0.1982594, 0.1982602, 0.1982598, 0.198261, 
    0.1982612, 0.1982615, 0.1982618, 0.1982618, 0.198262, 0.1982617, 
    0.198262, 0.1982609, 0.1982614, 0.1982601, 0.1982604, 0.1982603, 
    0.1982601, 0.1982606, 0.1982611, 0.1982611, 0.1982613, 0.1982618, 
    0.198261, 0.1982635, 0.1982619, 0.1982596, 0.1982601, 0.1982602, 0.19826, 
    0.1982612, 0.1982608, 0.198262, 0.1982617, 0.1982622, 0.1982619, 
    0.1982619, 0.1982615, 0.1982613, 0.1982608, 0.1982604, 0.19826, 
    0.1982601, 0.1982605, 0.1982612, 0.1982618, 0.1982617, 0.1982622, 
    0.1982609, 0.1982614, 0.1982612, 0.1982618, 0.1982606, 0.1982616, 
    0.1982603, 0.1982604, 0.1982608, 0.1982614, 0.1982616, 0.1982618, 
    0.1982617, 0.1982612, 0.1982611, 0.1982608, 0.1982607, 0.1982604, 
    0.1982602, 0.1982604, 0.1982606, 0.1982612, 0.1982617, 0.1982623, 
    0.1982625, 0.1982631, 0.1982626, 0.1982635, 0.1982627, 0.1982641, 
    0.1982616, 0.1982627, 0.1982608, 0.198261, 0.1982614, 0.1982622, 
    0.1982618, 0.1982623, 0.1982611, 0.1982605, 0.1982603, 0.19826, 
    0.1982603, 0.1982603, 0.1982606, 0.1982605, 0.1982612, 0.1982608, 
    0.1982619, 0.1982623, 0.1982634, 0.1982641, 0.1982648, 0.1982651, 
    0.1982652, 0.1982653,
  0.1985151, 0.1985151, 0.1985151, 0.1985152, 0.1985151, 0.1985152, 
    0.1985151, 0.1985151, 0.1985151, 0.1985151, 0.1985152, 0.1985152, 
    0.1985153, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985151, 0.1985151, 0.1985151, 0.1985151, 0.1985151, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985153, 0.1985152, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985152, 0.1985153, 
    0.1985152, 0.1985151, 0.1985151, 0.1985151, 0.1985151, 0.1985151, 
    0.1985151, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985152, 0.1985152, 0.1985152, 0.1985151, 0.1985151, 0.1985151, 
    0.1985151, 0.1985151, 0.1985152, 0.1985151, 0.1985152, 0.1985152, 
    0.1985153, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985153, 0.1985153, 0.1985151, 0.1985151, 0.1985152, 0.1985151, 
    0.1985151, 0.1985151, 0.1985151, 0.1985151, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985151, 0.1985151, 
    0.1985151, 0.1985151, 0.1985151, 0.1985151, 0.1985151, 0.1985152, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985151, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985153, 0.1985152, 0.1985153, 0.1985152, 0.1985152, 
    0.1985153, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985153, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985154, 0.1985154, 0.1985155, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985152, 0.1985153, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985155, 0.1985155, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985152, 0.1985153, 0.1985152, 0.1985152, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985153, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985152, 
    0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985153, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985152, 
    0.1985153, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985155, 0.1985155, 
    0.1985155, 0.1985155,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.609447, 8.609521, 8.609507, 8.609565, 8.609533, 8.609571, 8.609463, 
    8.609523, 8.609485, 8.609455, 8.609674, 8.609568, 8.609794, 8.609723, 
    8.609902, 8.609782, 8.609927, 8.6099, 8.609983, 8.60996, 8.610062, 
    8.609994, 8.610117, 8.610046, 8.610057, 8.609992, 8.609591, 8.609661, 
    8.609587, 8.609596, 8.609592, 8.609533, 8.609503, 8.609444, 8.609454, 
    8.609498, 8.609601, 8.609568, 8.609655, 8.609653, 8.609749, 8.609706, 
    8.609872, 8.609825, 8.609961, 8.609926, 8.609959, 8.609949, 8.609959, 
    8.609909, 8.60993, 8.609887, 8.609714, 8.609764, 8.609614, 8.609523, 
    8.609466, 8.609424, 8.609429, 8.609441, 8.609499, 8.609555, 8.609597, 
    8.609625, 8.609653, 8.609732, 8.609779, 8.60988, 8.609863, 8.609893, 
    8.609923, 8.609972, 8.609964, 8.609985, 8.609894, 8.609954, 8.609854, 
    8.609881, 8.609654, 8.609576, 8.609539, 8.609509, 8.609434, 8.609486, 
    8.609465, 8.609515, 8.609546, 8.609531, 8.609626, 8.609589, 8.609782, 
    8.609698, 8.60992, 8.609867, 8.609933, 8.6099, 8.609956, 8.609905, 
    8.609993, 8.610012, 8.609999, 8.61005, 8.609902, 8.609959, 8.60953, 
    8.609532, 8.609545, 8.609491, 8.609488, 8.609443, 8.609484, 8.609502, 
    8.609549, 8.609574, 8.6096, 8.609655, 8.609716, 8.609806, 8.609871, 
    8.609913, 8.609887, 8.60991, 8.609884, 8.609873, 8.610004, 8.60993, 
    8.610043, 8.610037, 8.609985, 8.610037, 8.609534, 8.60952, 8.609469, 
    8.609509, 8.609438, 8.609477, 8.609499, 8.609589, 8.60961, 8.609627, 
    8.609663, 8.609708, 8.609789, 8.60986, 8.609925, 8.609921, 8.609922, 
    8.609936, 8.6099, 8.609942, 8.609948, 8.609931, 8.610036, 8.610006, 
    8.610037, 8.610017, 8.609525, 8.60955, 8.609536, 8.60956, 8.609543, 
    8.609619, 8.609642, 8.60975, 8.609707, 8.609777, 8.609715, 8.609725, 
    8.609777, 8.609718, 8.609855, 8.609759, 8.609937, 8.60984, 8.609942, 
    8.609925, 8.609955, 8.609981, 8.610014, 8.610075, 8.610061, 8.610112, 
    8.609586, 8.609616, 8.609614, 8.609647, 8.609671, 8.609724, 8.60981, 
    8.609777, 8.609838, 8.609849, 8.609758, 8.609814, 8.609637, 8.609664, 
    8.609649, 8.609588, 8.609783, 8.609681, 8.609872, 8.609817, 8.609977, 
    8.609896, 8.610053, 8.610117, 8.610182, 8.610252, 8.609633, 8.609612, 
    8.609652, 8.609702, 8.609752, 8.609819, 8.609827, 8.609838, 8.609871, 
    8.609899, 8.609841, 8.609905, 8.609669, 8.609793, 8.609604, 8.609659, 
    8.609699, 8.609683, 8.609775, 8.609796, 8.609881, 8.609838, 8.610101, 
    8.609984, 8.610309, 8.610218, 8.609606, 8.609634, 8.609733, 8.609686, 
    8.609824, 8.609858, 8.609886, 8.609921, 8.609924, 8.609945, 8.609912, 
    8.609944, 8.609819, 8.609876, 8.609722, 8.609759, 8.609742, 8.609724, 
    8.609782, 8.609842, 8.609845, 8.609864, 8.609915, 8.609825, 8.610112, 
    8.609933, 8.609665, 8.609718, 8.609728, 8.609707, 8.609855, 8.609801, 
    8.609944, 8.609906, 8.60997, 8.609939, 8.609934, 8.609893, 8.609868, 
    8.609803, 8.60975, 8.60971, 8.609719, 8.609764, 8.609846, 8.609924, 
    8.609907, 8.609965, 8.609815, 8.609877, 8.609852, 8.609917, 8.609776, 
    8.609891, 8.609746, 8.609759, 8.6098, 8.609879, 8.6099, 8.609919, 
    8.609907, 8.609849, 8.609839, 8.609799, 8.609787, 8.609756, 8.609731, 
    8.609754, 8.609778, 8.609849, 8.609912, 8.609981, 8.609998, 8.610074, 
    8.61001, 8.610113, 8.610023, 8.610181, 8.6099, 8.610023, 8.609802, 
    8.609827, 8.609869, 8.609968, 8.609917, 8.609978, 8.609839, 8.609765, 
    8.609747, 8.609713, 8.609748, 8.609745, 8.60978, 8.609769, 8.609852, 
    8.609808, 8.609933, 8.609978, 8.610106, 8.610184, 8.610265, 8.610299, 
    8.610311, 8.610314 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  4.009688e-15, 4.010079e-15, 4.010008e-15, 4.010308e-15, 4.010145e-15, 
    4.010339e-15, 4.009768e-15, 4.010091e-15, 4.009882e-15, 4.009726e-15, 
    4.010881e-15, 4.010323e-15, 4.011498e-15, 4.011135e-15, 4.012059e-15, 
    4.011437e-15, 4.012186e-15, 4.012049e-15, 4.012481e-15, 4.012358e-15, 
    4.012894e-15, 4.012538e-15, 4.013185e-15, 4.012813e-15, 4.012868e-15, 
    4.012525e-15, 4.010443e-15, 4.010809e-15, 4.010419e-15, 4.010472e-15, 
    4.01045e-15, 4.010145e-15, 4.009986e-15, 4.009664e-15, 4.009721e-15, 
    4.009965e-15, 4.010496e-15, 4.010321e-15, 4.010778e-15, 4.010768e-15, 
    4.011272e-15, 4.011044e-15, 4.0119e-15, 4.011659e-15, 4.012363e-15, 
    4.012185e-15, 4.012353e-15, 4.012303e-15, 4.012354e-15, 4.012092e-15, 
    4.012204e-15, 4.011977e-15, 4.011086e-15, 4.011345e-15, 4.010568e-15, 
    4.010091e-15, 4.00978e-15, 4.009563e-15, 4.009594e-15, 4.00965e-15, 
    4.009966e-15, 4.010257e-15, 4.010476e-15, 4.010622e-15, 4.010766e-15, 
    4.011183e-15, 4.011423e-15, 4.011944e-15, 4.011857e-15, 4.012011e-15, 
    4.012167e-15, 4.01242e-15, 4.01238e-15, 4.01249e-15, 4.012011e-15, 
    4.012327e-15, 4.011806e-15, 4.011947e-15, 4.010778e-15, 4.010369e-15, 
    4.010172e-15, 4.01002e-15, 4.009617e-15, 4.009884e-15, 4.009778e-15, 
    4.010051e-15, 4.010211e-15, 4.010133e-15, 4.010626e-15, 4.010433e-15, 
    4.011437e-15, 4.011004e-15, 4.012149e-15, 4.011876e-15, 4.012215e-15, 
    4.012043e-15, 4.012336e-15, 4.012073e-15, 4.012533e-15, 4.012631e-15, 
    4.012563e-15, 4.01283e-15, 4.012057e-15, 4.012351e-15, 4.010129e-15, 
    4.010142e-15, 4.010204e-15, 4.009931e-15, 4.009902e-15, 4.009661e-15, 
    4.009878e-15, 4.009983e-15, 4.010222e-15, 4.010359e-15, 4.010491e-15, 
    4.010782e-15, 4.011102e-15, 4.01156e-15, 4.011893e-15, 4.012115e-15, 
    4.011981e-15, 4.012099e-15, 4.011966e-15, 4.011905e-15, 4.012592e-15, 
    4.012203e-15, 4.012792e-15, 4.01276e-15, 4.012492e-15, 4.012764e-15, 
    4.010151e-15, 4.010078e-15, 4.009801e-15, 4.010021e-15, 4.009635e-15, 
    4.00984e-15, 4.009969e-15, 4.010431e-15, 4.010539e-15, 4.010631e-15, 
    4.010818e-15, 4.011056e-15, 4.011472e-15, 4.011838e-15, 4.012177e-15, 
    4.012153e-15, 4.012161e-15, 4.012234e-15, 4.01205e-15, 4.012265e-15, 
    4.012298e-15, 4.012207e-15, 4.012756e-15, 4.012599e-15, 4.01276e-15, 
    4.012658e-15, 4.010103e-15, 4.010227e-15, 4.010159e-15, 4.010285e-15, 
    4.010194e-15, 4.010591e-15, 4.010709e-15, 4.011275e-15, 4.01105e-15, 
    4.011416e-15, 4.011089e-15, 4.011145e-15, 4.011416e-15, 4.011108e-15, 
    4.011813e-15, 4.011325e-15, 4.012237e-15, 4.011738e-15, 4.012268e-15, 
    4.012176e-15, 4.012331e-15, 4.012467e-15, 4.012643e-15, 4.01296e-15, 
    4.012888e-15, 4.013158e-15, 4.010416e-15, 4.010575e-15, 4.010566e-15, 
    4.010736e-15, 4.010861e-15, 4.011138e-15, 4.011579e-15, 4.011415e-15, 
    4.011721e-15, 4.011781e-15, 4.011319e-15, 4.011598e-15, 4.010685e-15, 
    4.010827e-15, 4.010746e-15, 4.010425e-15, 4.011446e-15, 4.010918e-15, 
    4.011897e-15, 4.011612e-15, 4.012446e-15, 4.012026e-15, 4.012847e-15, 
    4.013185e-15, 4.013528e-15, 4.013901e-15, 4.010667e-15, 4.010559e-15, 
    4.010758e-15, 4.011025e-15, 4.011288e-15, 4.011629e-15, 4.011667e-15, 
    4.011729e-15, 4.011897e-15, 4.012036e-15, 4.011744e-15, 4.012072e-15, 
    4.010849e-15, 4.011494e-15, 4.010513e-15, 4.010801e-15, 4.011011e-15, 
    4.010924e-15, 4.011398e-15, 4.011507e-15, 4.011952e-15, 4.011725e-15, 
    4.013096e-15, 4.012488e-15, 4.014203e-15, 4.013719e-15, 4.010519e-15, 
    4.010669e-15, 4.011185e-15, 4.01094e-15, 4.011654e-15, 4.011828e-15, 
    4.011974e-15, 4.012152e-15, 4.012175e-15, 4.012281e-15, 4.012106e-15, 
    4.012276e-15, 4.01163e-15, 4.011919e-15, 4.011132e-15, 4.011321e-15, 
    4.011235e-15, 4.011139e-15, 4.011438e-15, 4.011747e-15, 4.011762e-15, 
    4.01186e-15, 4.012121e-15, 4.011658e-15, 4.01316e-15, 4.012216e-15, 
    4.010833e-15, 4.011111e-15, 4.011161e-15, 4.011051e-15, 4.01181e-15, 
    4.011534e-15, 4.012279e-15, 4.01208e-15, 4.012409e-15, 4.012245e-15, 
    4.01222e-15, 4.012011e-15, 4.011878e-15, 4.011545e-15, 4.011277e-15, 
    4.011068e-15, 4.011117e-15, 4.011347e-15, 4.011768e-15, 4.012173e-15, 
    4.012083e-15, 4.012384e-15, 4.011603e-15, 4.011925e-15, 4.011798e-15, 
    4.012132e-15, 4.011409e-15, 4.012e-15, 4.011255e-15, 4.011322e-15, 
    4.011529e-15, 4.011942e-15, 4.012046e-15, 4.012142e-15, 4.012084e-15, 
    4.01178e-15, 4.011734e-15, 4.011526e-15, 4.011464e-15, 4.011308e-15, 
    4.011174e-15, 4.011294e-15, 4.011418e-15, 4.011784e-15, 4.012109e-15, 
    4.012467e-15, 4.012558e-15, 4.012956e-15, 4.01262e-15, 4.013163e-15, 
    4.012684e-15, 4.013523e-15, 4.012046e-15, 4.012687e-15, 4.011541e-15, 
    4.011666e-15, 4.011884e-15, 4.012402e-15, 4.012131e-15, 4.012452e-15, 
    4.011733e-15, 4.011351e-15, 4.011261e-15, 4.011079e-15, 4.011266e-15, 
    4.011251e-15, 4.011429e-15, 4.011373e-15, 4.011796e-15, 4.011569e-15, 
    4.012217e-15, 4.012452e-15, 4.013126e-15, 4.013536e-15, 4.013967e-15, 
    4.014153e-15, 4.01421e-15, 4.014234e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  11.11592, 11.16022, 11.1516, 11.1874, 11.16753, 11.19098, 11.12489, 
    11.16199, 11.1383, 11.1199, 11.25706, 11.18899, 11.32797, 11.28438, 
    11.39404, 11.32119, 11.40876, 11.39193, 11.44261, 11.42808, 11.49307, 
    11.44933, 11.52682, 11.48261, 11.48952, 11.44789, 11.20266, 11.24857, 
    11.19995, 11.20649, 11.20355, 11.16794, 11.15003, 11.11254, 11.11934, 
    11.14687, 11.20943, 11.18816, 11.24178, 11.24057, 11.30043, 11.27342, 
    11.3743, 11.34557, 11.42869, 11.40775, 11.4277, 11.42165, 11.42778, 
    11.39709, 11.41024, 11.38325, 11.27848, 11.30921, 11.21769, 11.16287, 
    11.12652, 11.10078, 11.10441, 11.11135, 11.14703, 11.18063, 11.20628, 
    11.22346, 11.24039, 11.29177, 11.319, 11.38012, 11.36907, 11.38779, 
    11.40567, 11.43575, 11.43079, 11.44406, 11.38729, 11.425, 11.36278, 
    11.37978, 11.24503, 11.1939, 11.17223, 11.15326, 11.10721, 11.139, 
    11.12646, 11.1563, 11.17528, 11.16589, 11.22393, 11.20134, 11.32062, 
    11.26915, 11.40359, 11.37133, 11.41132, 11.39091, 11.4259, 11.3944, 
    11.44899, 11.4609, 11.45276, 11.48403, 11.39266, 11.42771, 11.16563, 
    11.16716, 11.1743, 11.14295, 11.14104, 11.11235, 11.13787, 11.14875, 
    11.17638, 11.19275, 11.20832, 11.2426, 11.28096, 11.33472, 11.37342, 
    11.39941, 11.38347, 11.39754, 11.38181, 11.37444, 11.45644, 11.41036, 
    11.47953, 11.4757, 11.44437, 11.47613, 11.16824, 11.15942, 11.12887, 
    11.15277, 11.10923, 11.1336, 11.14762, 11.20182, 11.21374, 11.22481, 
    11.24669, 11.2748, 11.32421, 11.3673, 11.40671, 11.40382, 11.40484, 
    11.41366, 11.39183, 11.41724, 11.42151, 11.41035, 11.47519, 11.45664, 
    11.47562, 11.46354, 11.16229, 11.17712, 11.1691, 11.18418, 11.17356, 
    11.22084, 11.23504, 11.3016, 11.27425, 11.31779, 11.27866, 11.28559, 
    11.31922, 11.28078, 11.36493, 11.30785, 11.414, 11.35687, 11.41758, 
    11.40654, 11.42482, 11.44122, 11.46185, 11.49999, 11.49115, 11.52308, 
    11.19925, 11.21853, 11.21682, 11.23702, 11.25196, 11.28439, 11.33652, 
    11.3169, 11.35293, 11.36017, 11.30544, 11.33903, 11.23144, 11.24879, 
    11.23845, 11.20077, 11.32143, 11.25942, 11.37407, 11.34036, 11.43888, 
    11.38983, 11.48629, 11.52767, 11.56667, 11.61236, 11.22905, 11.21594, 
    11.23942, 11.27195, 11.30217, 11.34242, 11.34654, 11.35409, 11.37366, 
    11.39013, 11.35648, 11.39426, 11.25283, 11.32682, 11.211, 11.24581, 
    11.27003, 11.25939, 11.31466, 11.32771, 11.38082, 11.35334, 11.51746, 
    11.44469, 11.6472, 11.59042, 11.21137, 11.229, 11.29052, 11.26123, 
    11.3451, 11.3658, 11.38264, 11.4042, 11.40652, 11.41931, 11.39837, 
    11.41848, 11.3425, 11.37642, 11.28347, 11.30606, 11.29566, 11.28427, 
    11.31945, 11.35701, 11.35781, 11.36987, 11.40391, 11.34544, 11.52689, 
    11.41466, 11.24826, 11.28232, 11.28718, 11.27398, 11.36373, 11.33116, 
    11.41899, 11.39522, 11.43419, 11.41481, 11.41197, 11.38711, 11.37166, 
    11.33266, 11.30098, 11.27589, 11.28172, 11.30929, 11.35931, 11.40674, 
    11.39634, 11.43122, 11.33901, 11.37763, 11.3627, 11.40166, 11.31638, 
    11.389, 11.29786, 11.30583, 11.33052, 11.38026, 11.39127, 11.40304, 
    11.39577, 11.36058, 11.35482, 11.32991, 11.32305, 11.3041, 11.28843, 
    11.30275, 11.3178, 11.36059, 11.39924, 11.44145, 11.45179, 11.50127, 
    11.461, 11.52751, 11.47097, 11.56894, 11.39321, 11.46929, 11.33164, 
    11.34642, 11.3732, 11.43472, 11.40147, 11.44036, 11.35459, 11.31025, 
    11.29878, 11.27741, 11.29926, 11.29749, 11.31842, 11.31169, 11.36201, 
    11.33496, 11.4119, 11.44005, 11.51973, 11.56874, 11.61872, 11.64083, 
    11.64756, 11.65038 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  2.972005e-09, 2.937562e-09, 2.944186e-09, 2.916931e-09, 2.931978e-09, 
    2.914236e-09, 2.964948e-09, 2.936212e-09, 2.954482e-09, 2.968868e-09, 
    2.865673e-09, 2.915729e-09, 2.815761e-09, 2.846171e-09, 2.771188e-09, 
    2.820441e-09, 2.761498e-09, 2.772585e-09, 2.739533e-09, 2.748909e-09, 
    2.707608e-09, 2.735231e-09, 2.686764e-09, 2.714148e-09, 2.70982e-09, 
    2.736153e-09, 2.905496e-09, 2.871794e-09, 2.907521e-09, 2.902651e-09, 
    2.904835e-09, 2.931664e-09, 2.945402e-09, 2.974679e-09, 2.969314e-09, 
    2.947837e-09, 2.900468e-09, 2.91635e-09, 2.876712e-09, 2.877593e-09, 
    2.834877e-09, 2.853953e-09, 2.784317e-09, 2.803706e-09, 2.748516e-09, 
    2.762157e-09, 2.749152e-09, 2.753081e-09, 2.749101e-09, 2.769171e-09, 
    2.760531e-09, 2.778346e-09, 2.850357e-09, 2.828745e-09, 2.894357e-09, 
    2.935542e-09, 2.963673e-09, 2.984016e-09, 2.98112e-09, 2.975618e-09, 
    2.947713e-09, 2.92203e-09, 2.902803e-09, 2.890105e-09, 2.87772e-09, 
    2.840961e-09, 2.821951e-09, 2.780432e-09, 2.787823e-09, 2.775331e-09, 
    2.763523e-09, 2.743952e-09, 2.747152e-09, 2.738607e-09, 2.775661e-09, 
    2.750906e-09, 2.792053e-09, 2.780657e-09, 2.87436e-09, 2.912046e-09, 
    2.928404e-09, 2.942909e-09, 2.978898e-09, 2.953935e-09, 2.963717e-09, 
    2.940572e-09, 2.92608e-09, 2.933227e-09, 2.88976e-09, 2.906479e-09, 
    2.820834e-09, 2.856996e-09, 2.764894e-09, 2.786303e-09, 2.759819e-09, 
    2.773261e-09, 2.750321e-09, 2.770947e-09, 2.735444e-09, 2.727851e-09, 
    2.733034e-09, 2.713252e-09, 2.7721e-09, 2.749151e-09, 2.933427e-09, 
    2.932258e-09, 2.92683e-09, 2.95087e-09, 2.952356e-09, 2.974825e-09, 
    2.954814e-09, 2.946386e-09, 2.925246e-09, 2.912905e-09, 2.901286e-09, 
    2.876114e-09, 2.848594e-09, 2.811123e-09, 2.784903e-09, 2.767642e-09, 
    2.778197e-09, 2.768873e-09, 2.779301e-09, 2.78422e-09, 2.730689e-09, 
    2.76045e-09, 2.716077e-09, 2.718489e-09, 2.738404e-09, 2.718217e-09, 
    2.931439e-09, 2.938174e-09, 2.961837e-09, 2.943281e-09, 2.977297e-09, 
    2.958142e-09, 2.947257e-09, 2.906124e-09, 2.897268e-09, 2.889109e-09, 
    2.873152e-09, 2.852969e-09, 2.818348e-09, 2.789009e-09, 2.76284e-09, 
    2.764738e-09, 2.764069e-09, 2.758294e-09, 2.77265e-09, 2.755953e-09, 
    2.753172e-09, 2.760455e-09, 2.718813e-09, 2.730561e-09, 2.718541e-09, 
    2.726175e-09, 2.935981e-09, 2.924689e-09, 2.930778e-09, 2.919351e-09, 
    2.927389e-09, 2.892033e-09, 2.881625e-09, 2.834061e-09, 2.853363e-09, 
    2.82279e-09, 2.850223e-09, 2.845316e-09, 2.8218e-09, 2.848726e-09, 
    2.790606e-09, 2.829699e-09, 2.75807e-09, 2.796044e-09, 2.755729e-09, 
    2.762952e-09, 2.751019e-09, 2.740431e-09, 2.727247e-09, 2.703298e-09, 
    2.708801e-09, 2.689052e-09, 2.908042e-09, 2.893735e-09, 2.894991e-09, 
    2.880179e-09, 2.869338e-09, 2.846165e-09, 2.80989e-09, 2.823405e-09, 
    2.79871e-09, 2.793812e-09, 2.831377e-09, 2.808173e-09, 2.884253e-09, 
    2.871635e-09, 2.879134e-09, 2.906906e-09, 2.820274e-09, 2.86397e-09, 
    2.784474e-09, 2.807262e-09, 2.741935e-09, 2.773974e-09, 2.711841e-09, 
    2.686242e-09, 2.662667e-09, 2.635701e-09, 2.885999e-09, 2.895641e-09, 
    2.878431e-09, 2.855002e-09, 2.833664e-09, 2.805859e-09, 2.803052e-09, 
    2.797924e-09, 2.784746e-09, 2.773776e-09, 2.796305e-09, 2.771041e-09, 
    2.868721e-09, 2.816555e-09, 2.899304e-09, 2.873792e-09, 2.856372e-09, 
    2.863986e-09, 2.82496e-09, 2.81594e-09, 2.779963e-09, 2.798428e-09, 
    2.692506e-09, 2.738203e-09, 2.615596e-09, 2.648566e-09, 2.899027e-09, 
    2.886033e-09, 2.841839e-09, 2.862669e-09, 2.804027e-09, 2.790016e-09, 
    2.778747e-09, 2.76449e-09, 2.762963e-09, 2.754607e-09, 2.768331e-09, 
    2.755147e-09, 2.805801e-09, 2.7829e-09, 2.846814e-09, 2.830944e-09, 
    2.83822e-09, 2.84625e-09, 2.821636e-09, 2.795946e-09, 2.795407e-09, 
    2.787287e-09, 2.764689e-09, 2.803795e-09, 2.686728e-09, 2.757644e-09, 
    2.872016e-09, 2.847634e-09, 2.844196e-09, 2.853556e-09, 2.791413e-09, 
    2.813563e-09, 2.754811e-09, 2.770408e-09, 2.744959e-09, 2.757537e-09, 
    2.759398e-09, 2.775777e-09, 2.786087e-09, 2.812538e-09, 2.834495e-09, 
    2.852195e-09, 2.848057e-09, 2.828693e-09, 2.794393e-09, 2.762823e-09, 
    2.769667e-09, 2.746874e-09, 2.808185e-09, 2.782091e-09, 2.792108e-09, 
    2.766163e-09, 2.823765e-09, 2.774528e-09, 2.836677e-09, 2.8311e-09, 
    2.814007e-09, 2.780338e-09, 2.773022e-09, 2.765251e-09, 2.770041e-09, 
    2.793536e-09, 2.797431e-09, 2.814421e-09, 2.819152e-09, 2.832312e-09, 
    2.843314e-09, 2.833257e-09, 2.822783e-09, 2.793527e-09, 2.767756e-09, 
    2.74028e-09, 2.733654e-09, 2.702504e-09, 2.727793e-09, 2.686344e-09, 
    2.72148e-09, 2.661317e-09, 2.771742e-09, 2.722538e-09, 2.813237e-09, 
    2.80313e-09, 2.785057e-09, 2.744618e-09, 2.766284e-09, 2.740987e-09, 
    2.797584e-09, 2.828028e-09, 2.836037e-09, 2.851111e-09, 2.835694e-09, 
    2.836941e-09, 2.822354e-09, 2.827023e-09, 2.792568e-09, 2.810954e-09, 
    2.759444e-09, 2.741186e-09, 2.691105e-09, 2.661432e-09, 2.632e-09, 
    2.619242e-09, 2.615387e-09, 2.61378e-09 ;

 W_SCALAR =
  0.6401834, 0.64178, 0.6414698, 0.6427564, 0.6420428, 0.6428851, 0.6405072, 
    0.6418434, 0.6409906, 0.6403272, 0.6452497, 0.6428137, 0.647774, 
    0.6462244, 0.6501129, 0.6475331, 0.6506324, 0.6500384, 0.6518248, 
    0.6513133, 0.6535954, 0.6520607, 0.6547763, 0.653229, 0.6534713, 
    0.6520101, 0.6433042, 0.6449468, 0.6432068, 0.6434412, 0.643336, 
    0.6420576, 0.6414129, 0.6400612, 0.6403067, 0.6412994, 0.6435466, 
    0.6427841, 0.6447045, 0.6446611, 0.6467957, 0.6458337, 0.6494156, 
    0.6483986, 0.6513346, 0.650597, 0.6513, 0.6510869, 0.6513028, 0.6502208, 
    0.6506845, 0.6497318, 0.646014, 0.6471079, 0.6438424, 0.6418749, 
    0.6405659, 0.6396363, 0.6397678, 0.6400183, 0.6413051, 0.6425137, 
    0.6434339, 0.6440491, 0.6446549, 0.6464873, 0.6474556, 0.6496211, 
    0.6492305, 0.6498921, 0.6505235, 0.6515832, 0.6514089, 0.6518754, 
    0.6498745, 0.6512048, 0.6490079, 0.6496092, 0.6448202, 0.6429898, 
    0.6422115, 0.6415294, 0.6398688, 0.6410159, 0.6405638, 0.6416389, 
    0.6423215, 0.6419839, 0.6440659, 0.643257, 0.647513, 0.6456816, 
    0.6504499, 0.6493106, 0.6507228, 0.6500024, 0.6512365, 0.6501259, 
    0.652049, 0.6524674, 0.6521816, 0.6532791, 0.6500643, 0.6513001, 
    0.6419745, 0.6420296, 0.6422861, 0.6411582, 0.6410892, 0.6400545, 
    0.6409751, 0.641367, 0.642361, 0.6429487, 0.6435071, 0.6447338, 
    0.6461025, 0.6480136, 0.6493846, 0.6503026, 0.6497397, 0.6502367, 
    0.6496812, 0.6494206, 0.6523107, 0.6506888, 0.6531214, 0.6529869, 
    0.6518866, 0.653002, 0.6420682, 0.6417513, 0.6406505, 0.641512, 
    0.6399418, 0.640821, 0.6413264, 0.6432739, 0.6437013, 0.6440976, 
    0.6448798, 0.645883, 0.6476408, 0.649168, 0.6505603, 0.6504583, 
    0.6504942, 0.6508051, 0.650035, 0.6509315, 0.6510819, 0.6506886, 
    0.6529688, 0.6523179, 0.652984, 0.6525602, 0.6418543, 0.6423874, 
    0.6420994, 0.6426411, 0.6422595, 0.6439553, 0.6444632, 0.6468371, 
    0.6458633, 0.6474126, 0.6460207, 0.6462675, 0.6474633, 0.6460959, 
    0.649084, 0.6470592, 0.6508172, 0.6487985, 0.6509436, 0.6505542, 
    0.6511987, 0.6517756, 0.6525009, 0.653838, 0.6535285, 0.6546457, 
    0.6431818, 0.6438726, 0.6438117, 0.6445342, 0.6450682, 0.6462247, 
    0.6480775, 0.6473811, 0.6486591, 0.6489156, 0.6469737, 0.6481665, 
    0.6443346, 0.6449547, 0.6445854, 0.6432364, 0.6475418, 0.6453342, 
    0.6494072, 0.6482137, 0.6516933, 0.6499643, 0.6533581, 0.6548061, 
    0.6561666, 0.657755, 0.6442493, 0.6437802, 0.64462, 0.6457812, 0.6468573, 
    0.6482866, 0.6484327, 0.6487002, 0.6493928, 0.6499749, 0.6487849, 
    0.6501208, 0.6450986, 0.6477331, 0.6436028, 0.6448482, 0.6457127, 
    0.6453335, 0.6473014, 0.6477648, 0.649646, 0.6486739, 0.654449, 
    0.6518975, 0.6589624, 0.6569928, 0.6436162, 0.6442477, 0.6464429, 
    0.6453989, 0.6483819, 0.649115, 0.6497105, 0.6504716, 0.6505536, 
    0.6510043, 0.6502658, 0.650975, 0.6482896, 0.6494904, 0.6461921, 
    0.6469958, 0.6466261, 0.6462205, 0.6474718, 0.6488037, 0.648832, 
    0.6492587, 0.6504608, 0.6483939, 0.6547782, 0.65084, 0.6449358, 
    0.6461508, 0.646324, 0.6458536, 0.6490415, 0.6478875, 0.6509932, 
    0.6501547, 0.6515283, 0.6508459, 0.6507455, 0.6498684, 0.649322, 
    0.6479405, 0.6468151, 0.6459218, 0.6461295, 0.6471106, 0.6488851, 
    0.6505612, 0.6501942, 0.6514239, 0.6481658, 0.6495333, 0.649005, 
    0.6503819, 0.6473626, 0.6499347, 0.6467043, 0.6469879, 0.6478645, 
    0.6496261, 0.6500152, 0.6504308, 0.6501743, 0.6489301, 0.648726, 
    0.6478432, 0.6475994, 0.6469261, 0.6463685, 0.646878, 0.647413, 
    0.6489305, 0.6502964, 0.6517838, 0.6521475, 0.6538827, 0.6524706, 
    0.6548001, 0.6528203, 0.6562451, 0.6500833, 0.6527616, 0.6479043, 
    0.6484286, 0.6493764, 0.6515468, 0.6503754, 0.6517451, 0.648718, 
    0.6471445, 0.6467368, 0.6459762, 0.6467542, 0.6466909, 0.6474349, 
    0.6471959, 0.6489809, 0.6480224, 0.6507431, 0.6517343, 0.6545287, 
    0.6562384, 0.6579758, 0.658742, 0.6589751, 0.6590725,
  0.6386679, 0.6403095, 0.6399905, 0.6413135, 0.6405797, 0.6414458, 
    0.6390008, 0.6403747, 0.6394978, 0.6388156, 0.643877, 0.6413724, 
    0.6464723, 0.6448792, 0.6488768, 0.6462246, 0.6494108, 0.6488002, 
    0.6506366, 0.6501108, 0.6524569, 0.6508792, 0.6536708, 0.6520802, 
    0.6523293, 0.6508272, 0.6418767, 0.6435655, 0.6417766, 0.6420176, 
    0.6419094, 0.640595, 0.6399321, 0.6385422, 0.6387946, 0.6398153, 
    0.6421259, 0.6413419, 0.6433164, 0.6432719, 0.6454664, 0.6444775, 
    0.6481599, 0.6471144, 0.6501328, 0.6493744, 0.6500972, 0.6498781, 
    0.6501001, 0.6489877, 0.6494644, 0.6484851, 0.6446628, 0.6457875, 
    0.6424301, 0.6404071, 0.6390612, 0.6381053, 0.6382405, 0.6384981, 
    0.6398213, 0.6410639, 0.6420101, 0.6426426, 0.6432655, 0.6451494, 
    0.6461449, 0.6483712, 0.6479696, 0.6486498, 0.649299, 0.6503883, 
    0.6502091, 0.6506888, 0.6486318, 0.6499993, 0.6477408, 0.648359, 
    0.6434354, 0.6415535, 0.6407532, 0.6400518, 0.6383443, 0.6395238, 
    0.639059, 0.6401644, 0.6408663, 0.6405192, 0.6426599, 0.6418281, 
    0.6462039, 0.644321, 0.6492233, 0.648052, 0.6495038, 0.6487632, 
    0.6500319, 0.6488901, 0.6508672, 0.6512973, 0.6510034, 0.6521317, 
    0.6488268, 0.6500973, 0.6405095, 0.6405661, 0.6408299, 0.6396702, 
    0.6395992, 0.6385353, 0.639482, 0.6398849, 0.640907, 0.6415112, 
    0.6420853, 0.6433466, 0.6447538, 0.6467186, 0.648128, 0.6490718, 
    0.6484932, 0.6490041, 0.6484329, 0.6481651, 0.6511362, 0.6494689, 
    0.6519695, 0.6518313, 0.6507002, 0.6518468, 0.6406059, 0.64028, 
    0.6391481, 0.640034, 0.6384194, 0.6393235, 0.6398431, 0.6418456, 
    0.642285, 0.6426925, 0.6434967, 0.6445281, 0.6463353, 0.6479053, 
    0.6493367, 0.6492319, 0.6492688, 0.6495884, 0.6487967, 0.6497183, 
    0.649873, 0.6494686, 0.6518127, 0.6511436, 0.6518283, 0.6513926, 
    0.6403859, 0.6409341, 0.6406379, 0.6411949, 0.6408026, 0.6425462, 
    0.6430684, 0.6455091, 0.6445078, 0.6461007, 0.6446697, 0.6449234, 
    0.6461529, 0.644747, 0.647819, 0.6457374, 0.6496008, 0.6475255, 
    0.6497307, 0.6493305, 0.649993, 0.6505861, 0.6513317, 0.6527063, 
    0.6523881, 0.6535366, 0.6417509, 0.6424611, 0.6423985, 0.6431413, 
    0.6436903, 0.6448795, 0.6467842, 0.6460683, 0.6473822, 0.6476459, 
    0.6456495, 0.6468757, 0.6429362, 0.6435736, 0.643194, 0.641807, 
    0.6462335, 0.6439639, 0.6481513, 0.6469243, 0.6505015, 0.648724, 
    0.6522129, 0.6537014, 0.6550999, 0.6567327, 0.6428484, 0.6423661, 
    0.6432295, 0.6444235, 0.6455298, 0.6469992, 0.6471494, 0.6474245, 
    0.6481366, 0.648735, 0.6475115, 0.648885, 0.6437217, 0.6464302, 
    0.6421837, 0.6434642, 0.6443531, 0.6439631, 0.6459864, 0.6464628, 
    0.6483968, 0.6473974, 0.6533343, 0.6507115, 0.6579739, 0.6559492, 
    0.6421975, 0.6428468, 0.6451038, 0.6440304, 0.6470972, 0.6478509, 
    0.6484632, 0.6492456, 0.6493299, 0.6497931, 0.6490339, 0.6497631, 
    0.6470023, 0.6482369, 0.6448458, 0.6456722, 0.6452921, 0.6448751, 
    0.6461616, 0.6475309, 0.6475599, 0.6479986, 0.6492344, 0.6471096, 
    0.6536728, 0.6496243, 0.6435543, 0.6448034, 0.6449815, 0.6444979, 
    0.6477754, 0.6465889, 0.6497818, 0.6489197, 0.6503319, 0.6496304, 
    0.6495271, 0.6486254, 0.6480637, 0.6466433, 0.6454864, 0.644568, 
    0.6447816, 0.6457902, 0.6476145, 0.6493376, 0.6489604, 0.6502246, 
    0.6468751, 0.6482809, 0.6477378, 0.6491533, 0.6460493, 0.6486936, 
    0.6453725, 0.645664, 0.6465653, 0.6483763, 0.6487763, 0.6492036, 
    0.6489399, 0.6476607, 0.647451, 0.6465434, 0.6462928, 0.6456006, 
    0.6450272, 0.6455511, 0.6461011, 0.6476612, 0.6490655, 0.6505945, 
    0.6509684, 0.6527522, 0.6513005, 0.6536953, 0.65166, 0.6551806, 
    0.6488464, 0.6515998, 0.6466063, 0.6471452, 0.6481196, 0.6503509, 
    0.6491466, 0.6505548, 0.6474428, 0.645825, 0.6454059, 0.6446239, 
    0.6454238, 0.6453587, 0.6461237, 0.6458779, 0.647713, 0.6467276, 
    0.6495246, 0.6505436, 0.6534163, 0.6551738, 0.6569597, 0.6577473, 
    0.6579869, 0.6580871,
  0.6424645, 0.6441363, 0.6438113, 0.6451588, 0.6444114, 0.6452935, 
    0.6428035, 0.6442026, 0.6433095, 0.642615, 0.6477703, 0.6452188, 
    0.6504153, 0.6487916, 0.6528667, 0.6501628, 0.6534111, 0.6527885, 
    0.6546612, 0.654125, 0.6565179, 0.6549087, 0.6577564, 0.6561337, 
    0.6563877, 0.6548556, 0.6457325, 0.647453, 0.6456305, 0.645876, 
    0.6457658, 0.6444269, 0.6437519, 0.6423365, 0.6425935, 0.6436329, 
    0.6459864, 0.6451878, 0.6471993, 0.6471539, 0.6493901, 0.6483822, 
    0.6521356, 0.6510698, 0.6541474, 0.6533741, 0.6541111, 0.6538876, 
    0.654114, 0.6529797, 0.6534658, 0.6524672, 0.6485711, 0.6497173, 
    0.6462963, 0.6442356, 0.6428649, 0.6418916, 0.6420292, 0.6422916, 
    0.643639, 0.6449046, 0.6458684, 0.6465127, 0.6471473, 0.649067, 
    0.6500816, 0.6523511, 0.6519417, 0.6526352, 0.6532971, 0.654408, 
    0.6542252, 0.6547144, 0.6526167, 0.6540112, 0.6517084, 0.6523387, 
    0.6473204, 0.6454033, 0.6445881, 0.6438738, 0.6421351, 0.6433361, 
    0.6428627, 0.6439884, 0.6447033, 0.6443498, 0.6465303, 0.645683, 
    0.6501417, 0.6482229, 0.6532199, 0.6520257, 0.653506, 0.6527508, 
    0.6540446, 0.6528803, 0.6548964, 0.6553351, 0.6550353, 0.6561863, 
    0.6528157, 0.6541111, 0.6443399, 0.6443976, 0.6446662, 0.6434851, 
    0.6434128, 0.6423295, 0.6432934, 0.6437038, 0.6447448, 0.6453602, 
    0.645945, 0.64723, 0.6486639, 0.6506664, 0.6521032, 0.6530655, 0.6524755, 
    0.6529964, 0.652414, 0.652141, 0.6551708, 0.6534704, 0.6560208, 
    0.6558797, 0.6547261, 0.6558957, 0.6444381, 0.6441061, 0.6429535, 
    0.6438556, 0.6422114, 0.6431321, 0.6436613, 0.6457009, 0.6461484, 
    0.6465636, 0.6473829, 0.6484339, 0.6502756, 0.6518762, 0.6533356, 
    0.6532287, 0.6532663, 0.6535922, 0.6527849, 0.6537247, 0.6538824, 
    0.6534701, 0.6558609, 0.6551782, 0.6558768, 0.6554323, 0.644214, 
    0.6447724, 0.6444707, 0.645038, 0.6446384, 0.6464145, 0.6469465, 
    0.6494336, 0.6484132, 0.6500365, 0.6485782, 0.6488367, 0.6500897, 
    0.648657, 0.6517881, 0.6496662, 0.6536049, 0.651489, 0.6537374, 
    0.6533293, 0.6540049, 0.6546097, 0.6553701, 0.6567724, 0.6564478, 
    0.6576195, 0.6456043, 0.6463279, 0.6462641, 0.6470208, 0.6475803, 
    0.6487919, 0.6507333, 0.6500036, 0.6513429, 0.6516116, 0.6495767, 
    0.6508266, 0.6468118, 0.6474613, 0.6470745, 0.6456615, 0.6501719, 
    0.647859, 0.6521269, 0.6508761, 0.6545235, 0.6527109, 0.6562691, 
    0.6577877, 0.6592149, 0.6608814, 0.6467225, 0.646231, 0.6471108, 
    0.6483272, 0.6494547, 0.6509525, 0.6511055, 0.651386, 0.6521119, 
    0.652722, 0.6514747, 0.6528749, 0.6476122, 0.6503724, 0.6460453, 
    0.6473498, 0.6482555, 0.6478581, 0.64992, 0.6504056, 0.6523772, 
    0.6513583, 0.6574131, 0.6547376, 0.6621486, 0.6600817, 0.6460593, 
    0.6467207, 0.6490205, 0.6479267, 0.6510523, 0.6518207, 0.6524449, 
    0.6532426, 0.6533286, 0.653801, 0.6530268, 0.6537704, 0.6509556, 
    0.6522142, 0.6487577, 0.6495998, 0.6492124, 0.6487874, 0.6500986, 
    0.6514944, 0.651524, 0.6519713, 0.6532313, 0.6510649, 0.6577585, 
    0.6536288, 0.6474416, 0.6487144, 0.6488959, 0.648403, 0.6517437, 
    0.6505342, 0.6537895, 0.6529104, 0.6543504, 0.653635, 0.6535298, 
    0.6526103, 0.6520376, 0.6505897, 0.6494104, 0.6484745, 0.6486922, 
    0.6497201, 0.6515797, 0.6533365, 0.6529519, 0.654241, 0.6508259, 
    0.6522591, 0.6517054, 0.6531485, 0.6499842, 0.6526799, 0.6492944, 
    0.6495915, 0.6505101, 0.6523563, 0.6527641, 0.6531999, 0.652931, 
    0.6516268, 0.651413, 0.6504878, 0.6502323, 0.6495268, 0.6489425, 
    0.6494764, 0.6500369, 0.6516273, 0.6530591, 0.6546183, 0.6549996, 
    0.6568192, 0.6553384, 0.6577815, 0.6557051, 0.6592972, 0.6528356, 
    0.6556436, 0.6505519, 0.6511012, 0.6520946, 0.6543698, 0.6531418, 
    0.6545778, 0.6514046, 0.6497556, 0.6493284, 0.6485315, 0.6493466, 
    0.6492804, 0.65006, 0.6498095, 0.6516801, 0.6506756, 0.6535272, 
    0.6545664, 0.6574968, 0.6592903, 0.6611131, 0.6619172, 0.6621618, 
    0.6622641,
  0.6480104, 0.6497337, 0.6493987, 0.6507881, 0.6500174, 0.6509271, 
    0.6483598, 0.6498021, 0.6488814, 0.6481655, 0.6534824, 0.65085, 
    0.6562133, 0.6545366, 0.6587461, 0.6559525, 0.659309, 0.6586654, 
    0.6606014, 0.6600469, 0.6625221, 0.6608574, 0.6638039, 0.6621245, 
    0.6623874, 0.6608024, 0.6513798, 0.6531549, 0.6512747, 0.6515279, 
    0.6514142, 0.6500334, 0.6493374, 0.6478785, 0.6481434, 0.6492147, 
    0.6516417, 0.650818, 0.6528931, 0.6528462, 0.6551546, 0.6541141, 
    0.6579906, 0.6568894, 0.6600701, 0.6592706, 0.6600326, 0.6598015, 
    0.6600356, 0.6588629, 0.6593654, 0.6583332, 0.654309, 0.6554924, 
    0.6519614, 0.6498361, 0.6484231, 0.64742, 0.6475618, 0.6478322, 0.649221, 
    0.6505259, 0.65152, 0.6521847, 0.6528395, 0.6548209, 0.6558686, 
    0.6582133, 0.6577902, 0.6585068, 0.659191, 0.6603395, 0.6601505, 
    0.6606565, 0.6584878, 0.6599293, 0.6575491, 0.6582004, 0.6530181, 
    0.6510402, 0.6501996, 0.6494631, 0.6476709, 0.6489087, 0.6484209, 
    0.6495813, 0.6503184, 0.6499538, 0.6522029, 0.6513287, 0.6559308, 
    0.6539495, 0.6591113, 0.657877, 0.659407, 0.6586263, 0.6599638, 
    0.6587601, 0.6608446, 0.6612984, 0.6609883, 0.6621789, 0.6586934, 
    0.6600326, 0.6499436, 0.6500031, 0.6502801, 0.6490624, 0.6489878, 
    0.6478713, 0.6488647, 0.6492878, 0.6503611, 0.6509959, 0.651599, 
    0.6529248, 0.6544048, 0.6564726, 0.657957, 0.6589516, 0.6583418, 
    0.6588802, 0.6582783, 0.6579961, 0.6611284, 0.6593701, 0.6620077, 
    0.6618618, 0.6606685, 0.6618783, 0.6500449, 0.6497027, 0.6485143, 
    0.6494443, 0.6477496, 0.6486984, 0.6492439, 0.6513472, 0.6518089, 
    0.6522372, 0.6530826, 0.6541673, 0.656069, 0.6577225, 0.6592308, 
    0.6591203, 0.6591592, 0.6594961, 0.6586616, 0.6596331, 0.6597961, 
    0.6593698, 0.6618423, 0.6611362, 0.6618587, 0.661399, 0.6498139, 
    0.6503896, 0.6500785, 0.6506635, 0.6502514, 0.6520833, 0.6526323, 
    0.6551994, 0.654146, 0.6558221, 0.6543162, 0.6545832, 0.655877, 
    0.6543976, 0.6576315, 0.6554397, 0.6595092, 0.6573224, 0.6596462, 
    0.6592243, 0.6599227, 0.6605482, 0.6613346, 0.6627854, 0.6624495, 
    0.6636621, 0.6512476, 0.651994, 0.6519282, 0.6527089, 0.6532863, 
    0.654537, 0.6565418, 0.655788, 0.6571714, 0.6574491, 0.6553472, 
    0.6566381, 0.6524933, 0.6531635, 0.6527644, 0.6513066, 0.6559619, 
    0.6535739, 0.6579816, 0.6566892, 0.660459, 0.6585851, 0.6622646, 
    0.6638362, 0.6653138, 0.6670401, 0.6524011, 0.6518941, 0.6528018, 
    0.6540573, 0.6552212, 0.6567681, 0.6569263, 0.657216, 0.657966, 
    0.6585966, 0.6573077, 0.6587546, 0.6533192, 0.656169, 0.6517025, 
    0.6530484, 0.6539832, 0.653573, 0.6557018, 0.6562033, 0.6582403, 
    0.6571874, 0.6634485, 0.6606804, 0.6683533, 0.6662116, 0.6517169, 
    0.6523993, 0.6547729, 0.6536438, 0.6568713, 0.6576651, 0.6583102, 
    0.6591347, 0.6592236, 0.659712, 0.6589116, 0.6596803, 0.6567714, 
    0.6580718, 0.6545016, 0.6553711, 0.6549711, 0.6545323, 0.6558862, 
    0.657328, 0.6573586, 0.6578208, 0.659123, 0.6568843, 0.6638059, 0.659534, 
    0.6531432, 0.6544569, 0.6546443, 0.6541355, 0.6575856, 0.6563361, 0.6597, 
    0.6587913, 0.66028, 0.6595404, 0.6594316, 0.6584811, 0.6578893, 
    0.6563934, 0.6551756, 0.6542093, 0.654434, 0.6554953, 0.6574161, 
    0.6592317, 0.6588342, 0.6601669, 0.6566374, 0.6581181, 0.657546, 
    0.6590375, 0.655768, 0.658553, 0.6550557, 0.6553625, 0.6563113, 
    0.6582186, 0.6586401, 0.6590905, 0.6588126, 0.6574648, 0.6572438, 
    0.6562881, 0.6560243, 0.6552957, 0.6546924, 0.6552437, 0.6558225, 
    0.6574653, 0.658945, 0.6605571, 0.6609514, 0.6628339, 0.6613018, 
    0.6638297, 0.6616811, 0.6653991, 0.658714, 0.6616175, 0.6563544, 
    0.6569219, 0.6579482, 0.6603001, 0.6590304, 0.6605152, 0.6572352, 
    0.655532, 0.6550909, 0.6542681, 0.6551097, 0.6550412, 0.6558463, 
    0.6555876, 0.6575198, 0.6564821, 0.6594289, 0.6605034, 0.6635351, 
    0.6653919, 0.6672802, 0.6681135, 0.668367, 0.6684731,
  0.6561805, 0.6580046, 0.6576499, 0.6591215, 0.658305, 0.6592688, 0.6565502, 
    0.6580771, 0.6571023, 0.6563446, 0.6619784, 0.6591871, 0.6648781, 
    0.6630973, 0.6675715, 0.6646011, 0.6681705, 0.6674856, 0.6695469, 
    0.6689563, 0.671594, 0.6698195, 0.6729614, 0.6711701, 0.6714503, 
    0.669761, 0.6597486, 0.6616309, 0.6596372, 0.6599055, 0.659785, 0.658322, 
    0.657585, 0.656041, 0.6563212, 0.6574552, 0.6600262, 0.6591532, 
    0.6613531, 0.6613034, 0.6637534, 0.6626487, 0.6667677, 0.6655967, 
    0.668981, 0.6681297, 0.668941, 0.668695, 0.6689442, 0.6676958, 0.6682307, 
    0.6671322, 0.6628556, 0.6641123, 0.660365, 0.6581131, 0.6566172, 
    0.655556, 0.655706, 0.655992, 0.6574618, 0.6588438, 0.6598971, 0.6606019, 
    0.6612963, 0.6633991, 0.664512, 0.6670046, 0.6665545, 0.6673169, 
    0.668045, 0.6692679, 0.6690666, 0.6696054, 0.6672966, 0.6688311, 
    0.6662982, 0.6669909, 0.6614857, 0.6593887, 0.6584981, 0.6577181, 
    0.6558214, 0.6571312, 0.6566148, 0.6578432, 0.6586239, 0.6582378, 
    0.6606211, 0.6596945, 0.6645779, 0.662474, 0.6679601, 0.6666469, 
    0.6682749, 0.6674441, 0.6688677, 0.6675864, 0.6698059, 0.6702895, 
    0.6699591, 0.6712281, 0.6675155, 0.668941, 0.658227, 0.65829, 0.6585833, 
    0.6572939, 0.657215, 0.6560333, 0.6570847, 0.6575325, 0.6586691, 
    0.6593416, 0.659981, 0.6613868, 0.6629573, 0.6651537, 0.666732, 
    0.6677902, 0.6671413, 0.6677142, 0.6670738, 0.6667736, 0.6701083, 
    0.6682357, 0.6710455, 0.67089, 0.6696183, 0.6709075, 0.6583342, 
    0.6579717, 0.6567138, 0.6576983, 0.6559047, 0.6569086, 0.6574861, 
    0.659714, 0.6602034, 0.6606575, 0.6615542, 0.6627052, 0.6647249, 
    0.6664826, 0.6680874, 0.6679698, 0.6680112, 0.6683698, 0.6674816, 
    0.6685156, 0.6686893, 0.6682354, 0.6708692, 0.6701166, 0.6708867, 
    0.6703966, 0.6580896, 0.6586993, 0.6583698, 0.6589895, 0.658553, 
    0.6604944, 0.6610765, 0.663801, 0.6626826, 0.6644625, 0.6628633, 
    0.6631467, 0.6645208, 0.6629497, 0.6663858, 0.6640563, 0.6683837, 
    0.6660571, 0.6685296, 0.6680804, 0.668824, 0.6694901, 0.6703281, 
    0.6718748, 0.6715165, 0.6728101, 0.6596085, 0.6603996, 0.6603299, 
    0.6611578, 0.6617702, 0.6630976, 0.6652272, 0.6644263, 0.6658966, 
    0.6661919, 0.663958, 0.6653296, 0.6609291, 0.66164, 0.6612166, 0.6596709, 
    0.664611, 0.6620754, 0.6667581, 0.665384, 0.6693951, 0.6674002, 
    0.6713194, 0.6729959, 0.6745735, 0.6764184, 0.6608313, 0.6602937, 
    0.6612563, 0.6625884, 0.6638243, 0.6654678, 0.6656359, 0.6659439, 
    0.6667416, 0.6674124, 0.6660414, 0.6675806, 0.6618052, 0.6648311, 
    0.6600906, 0.6615179, 0.6625098, 0.6620745, 0.6643347, 0.6648676, 
    0.6670333, 0.6659136, 0.6725821, 0.669631, 0.6778231, 0.6755328, 
    0.6601059, 0.6608294, 0.6633481, 0.6621496, 0.6655775, 0.6664215, 
    0.6671077, 0.6679851, 0.6680797, 0.6685996, 0.6677477, 0.6685659, 
    0.6654713, 0.666854, 0.6630601, 0.6639834, 0.6635585, 0.6630927, 
    0.6645306, 0.666063, 0.6660956, 0.6665871, 0.6679726, 0.6655914, 
    0.6729636, 0.6684101, 0.6616185, 0.6630126, 0.6632115, 0.6626715, 
    0.666337, 0.6650086, 0.6685869, 0.6676196, 0.6692045, 0.6684169, 
    0.668301, 0.6672896, 0.66666, 0.6650695, 0.6637757, 0.6627498, 0.6629883, 
    0.6641153, 0.6661567, 0.6680884, 0.6676652, 0.6690841, 0.6653289, 
    0.6669034, 0.6662948, 0.6678816, 0.664405, 0.667366, 0.6636484, 
    0.6639743, 0.6649823, 0.6670103, 0.6674588, 0.667938, 0.6676422, 
    0.6662085, 0.6659736, 0.6649577, 0.6646773, 0.6639033, 0.6632627, 
    0.663848, 0.6644629, 0.666209, 0.6677831, 0.6694996, 0.6699197, 
    0.6719264, 0.6702931, 0.672989, 0.6706973, 0.6746646, 0.6675373, 
    0.6706295, 0.665028, 0.6656312, 0.6667226, 0.6692259, 0.6678742, 
    0.669455, 0.6659644, 0.6641543, 0.6636858, 0.6628122, 0.6637058, 
    0.663633, 0.6644883, 0.6642134, 0.666267, 0.6651638, 0.6682982, 
    0.6694424, 0.6726746, 0.6746569, 0.6766752, 0.6775665, 0.6778378, 
    0.6779513,
  0.6732582, 0.6752669, 0.674876, 0.6764984, 0.675598, 0.6766608, 0.673665, 
    0.6753467, 0.6742728, 0.6734388, 0.6796542, 0.6765708, 0.6828661, 
    0.6808925, 0.6858574, 0.6825588, 0.6865239, 0.6857619, 0.6880565, 
    0.6873986, 0.6903399, 0.6883603, 0.6918678, 0.6898666, 0.6901795, 
    0.6882951, 0.6771904, 0.6792699, 0.6770673, 0.6773636, 0.6772306, 
    0.6756167, 0.6748044, 0.6731048, 0.6734131, 0.6746615, 0.6774968, 
    0.6765333, 0.6789628, 0.6789079, 0.6816193, 0.6803959, 0.6849639, 
    0.6836634, 0.687426, 0.6864784, 0.6873815, 0.6871076, 0.6873851, 
    0.6859957, 0.6865907, 0.685369, 0.6806249, 0.6820169, 0.677871, 
    0.6753864, 0.6737388, 0.6725714, 0.6727363, 0.6730509, 0.6746688, 
    0.676192, 0.6773543, 0.6781326, 0.6788999, 0.6812268, 0.68246, 0.6852272, 
    0.6847271, 0.6855744, 0.6863842, 0.6877456, 0.6875214, 0.6881217, 
    0.6855518, 0.6872591, 0.6844423, 0.685212, 0.6791094, 0.6767932, 
    0.6758108, 0.6749511, 0.6728632, 0.6743047, 0.6737362, 0.675089, 
    0.6759496, 0.6755238, 0.6781539, 0.6771306, 0.6825331, 0.6802026, 
    0.6862897, 0.6848297, 0.68664, 0.6857157, 0.6872999, 0.685874, 0.6883452, 
    0.6888842, 0.6885158, 0.6899313, 0.6857951, 0.6873816, 0.675512, 
    0.6755814, 0.6759048, 0.6744838, 0.6743969, 0.6730963, 0.6742535, 
    0.6747467, 0.6759994, 0.6767412, 0.6774469, 0.679, 0.6807375, 0.6831718, 
    0.6849242, 0.6861007, 0.6853791, 0.6860162, 0.6853041, 0.6849704, 
    0.6886823, 0.6865963, 0.6897276, 0.6895541, 0.688136, 0.6895736, 
    0.6756301, 0.6752307, 0.6738452, 0.6749293, 0.6729547, 0.6740596, 
    0.6746955, 0.6771522, 0.6776925, 0.678194, 0.6791851, 0.6804585, 
    0.6826962, 0.6846471, 0.6864313, 0.6863005, 0.6863465, 0.6867456, 
    0.6857575, 0.6869079, 0.6871012, 0.686596, 0.6895308, 0.6886914, 
    0.6895504, 0.6890038, 0.6753604, 0.6760327, 0.6756694, 0.6763528, 
    0.6758714, 0.6780139, 0.6786571, 0.681672, 0.6804334, 0.6824052, 
    0.6806335, 0.6809472, 0.6824698, 0.6807291, 0.6845396, 0.6819549, 
    0.6867611, 0.6841745, 0.6869234, 0.6864236, 0.6872513, 0.6879932, 
    0.6889273, 0.6906534, 0.6902534, 0.6916987, 0.6770357, 0.6779092, 
    0.6778321, 0.6787469, 0.679424, 0.6808929, 0.6832533, 0.682365, 
    0.6839963, 0.6843242, 0.681846, 0.683367, 0.6784942, 0.67928, 0.6788119, 
    0.6771047, 0.6825699, 0.6797615, 0.6849533, 0.6834273, 0.6878874, 
    0.6856669, 0.6900333, 0.6919064, 0.693672, 0.6957404, 0.6783861, 
    0.6777923, 0.6788557, 0.6803291, 0.6816977, 0.6835204, 0.6837069, 
    0.6840489, 0.6849349, 0.6856806, 0.6841571, 0.6858675, 0.6794626, 
    0.6828139, 0.677568, 0.679145, 0.6802422, 0.6797606, 0.6822635, 
    0.6828544, 0.6852591, 0.6840152, 0.6914439, 0.6881502, 0.697318, 
    0.6947469, 0.6775849, 0.678384, 0.6811703, 0.6798437, 0.6836421, 
    0.6845793, 0.6853418, 0.6863175, 0.6864228, 0.6870014, 0.6860535, 
    0.6869639, 0.6835243, 0.6850598, 0.6808513, 0.6818741, 0.6814034, 
    0.6808875, 0.6824807, 0.6841812, 0.6842173, 0.6847632, 0.6863036, 
    0.6836575, 0.6918702, 0.6867904, 0.6792561, 0.6807988, 0.6810191, 
    0.6804211, 0.6844853, 0.6830108, 0.6869873, 0.6859109, 0.6876751, 
    0.686798, 0.6866691, 0.685544, 0.6848442, 0.6830785, 0.681644, 0.6805078, 
    0.6807718, 0.6820203, 0.6842852, 0.6864324, 0.6859617, 0.6875408, 
    0.6833662, 0.6851147, 0.6844386, 0.6862023, 0.6823415, 0.685629, 
    0.681503, 0.681864, 0.6829816, 0.6852335, 0.6857321, 0.6862651, 
    0.6859362, 0.6843427, 0.6840818, 0.6829544, 0.6826434, 0.6817853, 
    0.6810756, 0.6817241, 0.6824057, 0.6843433, 0.6860929, 0.6880038, 
    0.6884719, 0.6907112, 0.6888883, 0.6918986, 0.6893391, 0.693774, 
    0.6858195, 0.6892635, 0.6830324, 0.6837018, 0.6849138, 0.6876988, 
    0.6861941, 0.687954, 0.6840715, 0.6820635, 0.6815444, 0.6805769, 
    0.6815665, 0.681486, 0.6824337, 0.682129, 0.6844077, 0.683183, 0.686666, 
    0.6879401, 0.6915472, 0.6937655, 0.6960286, 0.6970297, 0.6973346, 
    0.6974621,
  0.6968738, 0.6993591, 0.6988748, 0.7008876, 0.6997698, 0.7010895, 
    0.6973764, 0.6994581, 0.698128, 0.6970968, 0.7048212, 0.7009776, 0.70885, 
    0.7063712, 0.7126261, 0.7084634, 0.7134706, 0.7125052, 0.7154173, 
    0.7145808, 0.7183295, 0.7158039, 0.7202864, 0.7177247, 0.7181244, 
    0.7157209, 0.7017481, 0.7043408, 0.701595, 0.7019636, 0.7017981, 
    0.6997929, 0.6987861, 0.6966842, 0.6970651, 0.6986091, 0.7021295, 
    0.7009311, 0.7039573, 0.7038887, 0.707283, 0.7057492, 0.7114957, 
    0.7098542, 0.7146157, 0.713413, 0.7145591, 0.7142112, 0.7145637, 
    0.7128012, 0.7135555, 0.7120079, 0.706036, 0.7077823, 0.7025955, 
    0.6995074, 0.6974676, 0.696026, 0.6962296, 0.6966178, 0.6986181, 
    0.700507, 0.7019521, 0.7029215, 0.7038788, 0.7067904, 0.7083392, 
    0.7118286, 0.7111964, 0.7122678, 0.7132936, 0.7150219, 0.7147369, 
    0.7155003, 0.7122393, 0.7144037, 0.7108368, 0.7118093, 0.7041403, 
    0.701254, 0.7000338, 0.6989679, 0.6963861, 0.6981674, 0.6974644, 
    0.6991387, 0.700206, 0.6996778, 0.702948, 0.7016737, 0.7084312, 
    0.7055072, 0.7131737, 0.7113261, 0.7136179, 0.7124467, 0.7144555, 
    0.7126472, 0.7157847, 0.7164713, 0.716002, 0.7178074, 0.7125472, 
    0.7145593, 0.699663, 0.6997491, 0.7001504, 0.6983892, 0.6982816, 
    0.6966739, 0.698104, 0.6987146, 0.7002679, 0.7011895, 0.7020673, 
    0.7040038, 0.7061771, 0.7092348, 0.7114456, 0.7129343, 0.7120208, 
    0.7128271, 0.7119258, 0.711504, 0.7162139, 0.7135625, 0.7175472, 
    0.7173256, 0.7155185, 0.7173506, 0.6998096, 0.6993142, 0.6975991, 
    0.6989408, 0.6964991, 0.6978643, 0.6986512, 0.7017005, 0.7023731, 
    0.7029981, 0.7042349, 0.7058275, 0.7086362, 0.7110954, 0.7133532, 
    0.7131873, 0.7132457, 0.7137519, 0.7124996, 0.7139578, 0.7142031, 
    0.7135621, 0.717296, 0.7162256, 0.7173209, 0.7166237, 0.6994752, 
    0.7003093, 0.6998584, 0.7007067, 0.7001089, 0.7027735, 0.7035757, 
    0.7073491, 0.7057962, 0.7082702, 0.7060468, 0.7064399, 0.7083516, 
    0.7061666, 0.7109596, 0.7077044, 0.7137715, 0.7104988, 0.7139775, 
    0.7133434, 0.7143937, 0.7153367, 0.7165262, 0.7187305, 0.7182189, 
    0.7200694, 0.7015556, 0.7026431, 0.7025471, 0.7036878, 0.7045333, 
    0.7063718, 0.7093375, 0.7082198, 0.710274, 0.7106877, 0.7075676, 
    0.7094806, 0.7033724, 0.7043534, 0.7037689, 0.7016414, 0.7084773, 
    0.7049553, 0.7114823, 0.7095567, 0.7152022, 0.7123849, 0.7179376, 
    0.7203358, 0.7226056, 0.7252764, 0.7032377, 0.7024974, 0.7038236, 
    0.7056656, 0.7073814, 0.7096739, 0.7099091, 0.7103403, 0.711459, 
    0.7124022, 0.7104769, 0.712639, 0.7045816, 0.7087843, 0.702218, 
    0.7041848, 0.7055567, 0.7049541, 0.7080922, 0.7088352, 0.7118689, 
    0.7102978, 0.7197427, 0.7155365, 0.7273219, 0.723992, 0.7022391, 
    0.703235, 0.7067197, 0.705058, 0.7098273, 0.7110098, 0.7119735, 0.713209, 
    0.7133424, 0.7140765, 0.7128744, 0.7140288, 0.7096788, 0.711617, 
    0.7063197, 0.7076029, 0.707012, 0.706365, 0.7083652, 0.7105072, 
    0.7105528, 0.7112421, 0.7131913, 0.7098467, 0.7202895, 0.7138087, 
    0.7043236, 0.7062539, 0.70653, 0.7057807, 0.7108911, 0.7090322, 
    0.7140585, 0.7126939, 0.7149322, 0.7138184, 0.7136548, 0.7122293, 
    0.7113444, 0.7091173, 0.7073139, 0.7058893, 0.7062201, 0.7077865, 
    0.7106385, 0.7133546, 0.7127581, 0.7147616, 0.7094796, 0.7116863, 
    0.7108321, 0.7130631, 0.7081901, 0.7123369, 0.707137, 0.7075902, 
    0.7089953, 0.7118366, 0.7124674, 0.7131426, 0.7127258, 0.7107111, 
    0.7103818, 0.7089611, 0.7085698, 0.7074915, 0.706601, 0.7074146, 
    0.7082708, 0.7107118, 0.7129243, 0.7153502, 0.7159461, 0.7188044, 
    0.7164764, 0.7203259, 0.7170513, 0.7227371, 0.7125781, 0.7169549, 
    0.7090593, 0.7099025, 0.7114323, 0.7149624, 0.7130526, 0.7152869, 
    0.7103689, 0.7078408, 0.7071889, 0.7059758, 0.7072167, 0.7071156, 
    0.7083061, 0.7079232, 0.7107931, 0.709249, 0.7136508, 0.7152691, 
    0.7198752, 0.722726, 0.7256495, 0.7269474, 0.7273434, 0.727509,
  0.7536336, 0.7576361, 0.7568524, 0.7601215, 0.7583021, 0.7604513, 
    0.7544393, 0.7577966, 0.7556475, 0.7539908, 0.7666051, 0.7602684, 
    0.7733832, 0.769196, 0.7798715, 0.7727266, 0.7813413, 0.7796615, 
    0.7847567, 0.7832844, 0.7899396, 0.7854396, 0.7934738, 0.7888559, 
    0.7895718, 0.7852929, 0.7615288, 0.7658064, 0.7612781, 0.7618824, 
    0.7616109, 0.7583396, 0.7567091, 0.7533303, 0.7539399, 0.7564232, 
    0.7621546, 0.7601925, 0.7651701, 0.7650564, 0.7707297, 0.7681537, 
    0.7779149, 0.7750956, 0.7833456, 0.7812408, 0.7832464, 0.7826362, 
    0.7832543, 0.7801757, 0.7814893, 0.7788, 0.7686339, 0.7715728, 0.7629209, 
    0.7578763, 0.7545856, 0.752279, 0.7526037, 0.753224, 0.7564378, 
    0.7595009, 0.7618635, 0.763458, 0.7650401, 0.7699003, 0.7725158, 
    0.7784898, 0.7773989, 0.7792498, 0.7810325, 0.7840599, 0.7835586, 
    0.7849032, 0.7792005, 0.7829735, 0.7767802, 0.7784564, 0.7654737, 
    0.7607201, 0.7587309, 0.7570028, 0.7528537, 0.7557111, 0.7545804, 
    0.7572792, 0.7590109, 0.7581527, 0.7635017, 0.7614071, 0.7726718, 
    0.7677492, 0.7808238, 0.7776223, 0.7815983, 0.7795601, 0.7830645, 
    0.779908, 0.7854056, 0.7866221, 0.7857901, 0.7890038, 0.7797344, 
    0.7832465, 0.7581288, 0.7582685, 0.7589206, 0.7560683, 0.755895, 
    0.7533137, 0.755609, 0.7565935, 0.7591116, 0.7606146, 0.7620526, 
    0.7652471, 0.7688702, 0.7740384, 0.7778285, 0.780407, 0.7788221, 
    0.7802207, 0.7786579, 0.7779292, 0.7861656, 0.7815017, 0.7885385, 
    0.7881429, 0.7849354, 0.7881874, 0.7583667, 0.7575634, 0.7547967, 
    0.756959, 0.7530343, 0.755223, 0.7564912, 0.761451, 0.7625551, 0.7635843, 
    0.7656305, 0.7682848, 0.7730199, 0.777225, 0.7811366, 0.7808475, 
    0.7809492, 0.7818323, 0.7796518, 0.7821925, 0.782622, 0.7815009, 
    0.7880899, 0.7861864, 0.7881345, 0.7868928, 0.7578242, 0.7591789, 
    0.7584459, 0.7598264, 0.758853, 0.7632141, 0.7645382, 0.7708413, 
    0.7682323, 0.7723989, 0.7686518, 0.7693112, 0.7725368, 0.7688526, 
    0.7769913, 0.7714411, 0.7818667, 0.7761997, 0.7822269, 0.7811195, 
    0.7829561, 0.7846147, 0.7867196, 0.7906604, 0.7897412, 0.7930799, 
    0.7612137, 0.7629992, 0.7628412, 0.7647237, 0.7661263, 0.7691969, 
    0.7742134, 0.7723134, 0.7758141, 0.7765239, 0.77121, 0.7744575, 
    0.7642021, 0.7658274, 0.764858, 0.7613541, 0.7727501, 0.7668285, 
    0.7778917, 0.7745873, 0.7843774, 0.7794529, 0.789237, 0.7935637, 
    0.7977186, 0.8026853, 0.7639796, 0.7627594, 0.7649485, 0.7680139, 
    0.7708958, 0.7747874, 0.7751894, 0.7759277, 0.7778516, 0.7794829, 
    0.776162, 0.7798937, 0.7662065, 0.7732716, 0.7623001, 0.7655474, 
    0.7678319, 0.7668266, 0.7720972, 0.7733582, 0.7785594, 0.7758549, 
    0.7924877, 0.7849671, 0.8065489, 0.800286, 0.7623347, 0.7639752, 
    0.7697812, 0.7669997, 0.7750496, 0.7770777, 0.7787403, 0.7808851, 
    0.7811177, 0.7824001, 0.7803028, 0.7823168, 0.7747958, 0.7781242, 
    0.7691095, 0.7712696, 0.7702731, 0.7691855, 0.7725599, 0.7762139, 
    0.7762922, 0.7774776, 0.7808545, 0.7750828, 0.7934794, 0.7819317, 
    0.7657779, 0.768999, 0.7694624, 0.7682065, 0.7768735, 0.7736932, 
    0.7823687, 0.7799891, 0.783902, 0.7819487, 0.7816628, 0.7791833, 
    0.7776541, 0.7738381, 0.7707819, 0.7683882, 0.7689424, 0.77158, 
    0.7764394, 0.7811391, 0.7801008, 0.7836021, 0.7744558, 0.7782439, 
    0.776772, 0.7806311, 0.7722632, 0.7793697, 0.7704836, 0.7712482, 
    0.7736306, 0.7785036, 0.779596, 0.7807695, 0.7800446, 0.7765641, 
    0.775999, 0.7735722, 0.7729072, 0.7710815, 0.7695817, 0.7709517, 
    0.7723999, 0.7765653, 0.7803896, 0.7846385, 0.7856911, 0.7907935, 
    0.7866313, 0.7935457, 0.7876538, 0.797961, 0.779788, 0.787482, 0.7737394, 
    0.7751782, 0.7778056, 0.7839553, 0.7806128, 0.7845268, 0.7759768, 
    0.7716718, 0.7705711, 0.7685331, 0.7706179, 0.7704476, 0.7724597, 
    0.7718111, 0.776705, 0.7740625, 0.7816558, 0.7844955, 0.7927276, 
    0.7979407, 0.8033861, 0.8058377, 0.8065898, 0.806905,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.698417e-11, 3.713944e-11, 3.710917e-11, 3.723446e-11, 3.716493e-11, 
    3.724689e-11, 3.701546e-11, 3.714531e-11, 3.706237e-11, 3.699784e-11, 
    3.747741e-11, 3.723975e-11, 3.772486e-11, 3.757293e-11, 3.795468e-11, 
    3.770108e-11, 3.800583e-11, 3.794733e-11, 3.812342e-11, 3.80729e-11, 
    3.829812e-11, 3.814661e-11, 3.841502e-11, 3.826189e-11, 3.828576e-11, 
    3.814141e-11, 3.728789e-11, 3.744808e-11, 3.727831e-11, 3.730116e-11, 
    3.729087e-11, 3.716617e-11, 3.710333e-11, 3.697198e-11, 3.699577e-11, 
    3.709224e-11, 3.731114e-11, 3.723677e-11, 3.742419e-11, 3.741996e-11, 
    3.762875e-11, 3.753455e-11, 3.788598e-11, 3.778597e-11, 3.807496e-11, 
    3.800217e-11, 3.807145e-11, 3.805038e-11, 3.807161e-11, 3.796497e-11, 
    3.801056e-11, 3.791677e-11, 3.755265e-11, 3.765977e-11, 3.734025e-11, 
    3.714824e-11, 3.702098e-11, 3.693073e-11, 3.69434e-11, 3.696772e-11, 
    3.709272e-11, 3.721038e-11, 3.730011e-11, 3.736009e-11, 3.741923e-11, 
    3.759836e-11, 3.769333e-11, 3.790607e-11, 3.786769e-11, 3.793267e-11, 
    3.799489e-11, 3.809928e-11, 3.808208e-11, 3.812804e-11, 3.793078e-11, 
    3.806181e-11, 3.784548e-11, 3.79046e-11, 3.743551e-11, 3.7257e-11, 
    3.7181e-11, 3.711462e-11, 3.695317e-11, 3.706462e-11, 3.702062e-11, 
    3.712516e-11, 3.719161e-11, 3.715868e-11, 3.736169e-11, 3.728266e-11, 
    3.76989e-11, 3.751948e-11, 3.798768e-11, 3.787548e-11, 3.801446e-11, 
    3.794352e-11, 3.8065e-11, 3.79556e-11, 3.814511e-11, 3.81864e-11, 
    3.815809e-11, 3.826658e-11, 3.794929e-11, 3.807103e-11, 3.715799e-11, 
    3.716335e-11, 3.718829e-11, 3.707839e-11, 3.707167e-11, 3.697108e-11, 
    3.70605e-11, 3.70986e-11, 3.719538e-11, 3.725257e-11, 3.730698e-11, 
    3.74268e-11, 3.75606e-11, 3.774794e-11, 3.78827e-11, 3.797302e-11, 
    3.791759e-11, 3.796645e-11, 3.791174e-11, 3.788606e-11, 3.817079e-11, 
    3.801082e-11, 3.825086e-11, 3.823758e-11, 3.812881e-11, 3.823896e-11, 
    3.716704e-11, 3.713613e-11, 3.702901e-11, 3.711276e-11, 3.696006e-11, 
    3.704547e-11, 3.709453e-11, 3.728421e-11, 3.732593e-11, 3.73646e-11, 
    3.7441e-11, 3.753907e-11, 3.771131e-11, 3.786128e-11, 3.799836e-11, 
    3.798825e-11, 3.799177e-11, 3.802232e-11, 3.794645e-11, 3.80347e-11, 
    3.804945e-11, 3.801072e-11, 3.823569e-11, 3.817138e-11, 3.823714e-11, 
    3.81952e-11, 3.714612e-11, 3.719797e-11, 3.716986e-11, 3.722262e-11, 
    3.718536e-11, 3.73507e-11, 3.740024e-11, 3.76325e-11, 3.753712e-11, 
    3.768893e-11, 3.755248e-11, 3.757663e-11, 3.769366e-11, 3.755975e-11, 
    3.785284e-11, 3.765393e-11, 3.802347e-11, 3.782458e-11, 3.803585e-11, 
    3.799744e-11, 3.806091e-11, 3.811779e-11, 3.818933e-11, 3.832149e-11, 
    3.82908e-11, 3.840141e-11, 3.727537e-11, 3.734267e-11, 3.733676e-11, 
    3.740725e-11, 3.745939e-11, 3.75726e-11, 3.775422e-11, 3.768584e-11, 
    3.781128e-11, 3.783647e-11, 3.764577e-11, 3.776275e-11, 3.738739e-11, 
    3.744787e-11, 3.741184e-11, 3.728005e-11, 3.770119e-11, 3.748484e-11, 
    3.788444e-11, 3.776708e-11, 3.810956e-11, 3.793911e-11, 3.827392e-11, 
    3.841715e-11, 3.855218e-11, 3.870983e-11, 3.737945e-11, 3.73336e-11, 
    3.741558e-11, 3.752907e-11, 3.763445e-11, 3.77747e-11, 3.778903e-11, 
    3.781524e-11, 3.788331e-11, 3.79406e-11, 3.782341e-11, 3.795485e-11, 
    3.746179e-11, 3.771998e-11, 3.731573e-11, 3.74373e-11, 3.752184e-11, 
    3.748476e-11, 3.767753e-11, 3.772292e-11, 3.790768e-11, 3.781216e-11, 
    3.838164e-11, 3.812946e-11, 3.883006e-11, 3.863401e-11, 3.731754e-11, 
    3.737914e-11, 3.759378e-11, 3.749161e-11, 3.778398e-11, 3.785602e-11, 
    3.791455e-11, 3.798944e-11, 3.799747e-11, 3.804186e-11, 3.796904e-11, 
    3.803893e-11, 3.777457e-11, 3.789264e-11, 3.756884e-11, 3.764751e-11, 
    3.761128e-11, 3.757148e-11, 3.769409e-11, 3.78248e-11, 3.782761e-11, 
    3.786946e-11, 3.798748e-11, 3.778443e-11, 3.841393e-11, 3.802475e-11, 
    3.744635e-11, 3.756506e-11, 3.758206e-11, 3.753603e-11, 3.784868e-11, 
    3.773531e-11, 3.804079e-11, 3.795812e-11, 3.809346e-11, 3.802617e-11, 
    3.801618e-11, 3.792982e-11, 3.787595e-11, 3.774018e-11, 3.762969e-11, 
    3.754225e-11, 3.75625e-11, 3.765859e-11, 3.78327e-11, 3.799768e-11, 
    3.796147e-11, 3.808266e-11, 3.776194e-11, 3.789631e-11, 3.784426e-11, 
    3.797981e-11, 3.768385e-11, 3.793636e-11, 3.761929e-11, 3.764702e-11, 
    3.773294e-11, 3.790599e-11, 3.79443e-11, 3.798521e-11, 3.79599e-11, 
    3.783743e-11, 3.781735e-11, 3.773061e-11, 3.770659e-11, 3.764061e-11, 
    3.758587e-11, 3.76358e-11, 3.768813e-11, 3.783719e-11, 3.797153e-11, 
    3.81181e-11, 3.815401e-11, 3.832527e-11, 3.818569e-11, 3.841589e-11, 
    3.821994e-11, 3.855923e-11, 3.795098e-11, 3.821514e-11, 3.773689e-11, 
    3.77883e-11, 3.788136e-11, 3.809508e-11, 3.797966e-11, 3.811463e-11, 
    3.781654e-11, 3.766194e-11, 3.762201e-11, 3.75475e-11, 3.762363e-11, 
    3.761744e-11, 3.769036e-11, 3.766685e-11, 3.784203e-11, 3.77479e-11, 
    3.801538e-11, 3.811311e-11, 3.838934e-11, 3.855877e-11, 3.873154e-11, 
    3.880776e-11, 3.883097e-11, 3.884063e-11,
  2.48181e-11, 2.494881e-11, 2.49234e-11, 2.502892e-11, 2.497039e-11, 
    2.503949e-11, 2.484461e-11, 2.495399e-11, 2.488416e-11, 2.482989e-11, 
    2.523398e-11, 2.503363e-11, 2.544277e-11, 2.531461e-11, 2.563694e-11, 
    2.542279e-11, 2.568018e-11, 2.56308e-11, 2.577963e-11, 2.573697e-11, 
    2.592748e-11, 2.579932e-11, 2.602645e-11, 2.589688e-11, 2.591712e-11, 
    2.579509e-11, 2.507396e-11, 2.5209e-11, 2.506596e-11, 2.50852e-11, 
    2.507657e-11, 2.497158e-11, 2.491868e-11, 2.480815e-11, 2.482821e-11, 
    2.490942e-11, 2.509386e-11, 2.503124e-11, 2.518923e-11, 2.518566e-11, 
    2.536184e-11, 2.528236e-11, 2.557902e-11, 2.549462e-11, 2.573875e-11, 
    2.567729e-11, 2.573586e-11, 2.57181e-11, 2.573609e-11, 2.564597e-11, 
    2.568457e-11, 2.560532e-11, 2.529723e-11, 2.538766e-11, 2.511821e-11, 
    2.495651e-11, 2.484939e-11, 2.477342e-11, 2.478416e-11, 2.480462e-11, 
    2.49099e-11, 2.500903e-11, 2.508464e-11, 2.513525e-11, 2.518515e-11, 
    2.533622e-11, 2.54164e-11, 2.559607e-11, 2.556366e-11, 2.56186e-11, 
    2.567118e-11, 2.575946e-11, 2.574493e-11, 2.578384e-11, 2.561719e-11, 
    2.572789e-11, 2.55452e-11, 2.559513e-11, 2.519855e-11, 2.504814e-11, 
    2.498414e-11, 2.492828e-11, 2.479241e-11, 2.488621e-11, 2.484921e-11, 
    2.493728e-11, 2.499326e-11, 2.496557e-11, 2.513664e-11, 2.507009e-11, 
    2.542115e-11, 2.526977e-11, 2.566505e-11, 2.557032e-11, 2.568777e-11, 
    2.562783e-11, 2.573055e-11, 2.56381e-11, 2.579833e-11, 2.583324e-11, 
    2.580938e-11, 2.590112e-11, 2.563297e-11, 2.573584e-11, 2.496479e-11, 
    2.49693e-11, 2.499035e-11, 2.489786e-11, 2.489221e-11, 2.480759e-11, 
    2.48829e-11, 2.491497e-11, 2.499652e-11, 2.504476e-11, 2.509065e-11, 
    2.519163e-11, 2.530452e-11, 2.546265e-11, 2.557645e-11, 2.56528e-11, 
    2.560599e-11, 2.564732e-11, 2.560111e-11, 2.557947e-11, 2.582014e-11, 
    2.568492e-11, 2.588792e-11, 2.587668e-11, 2.578475e-11, 2.587795e-11, 
    2.497248e-11, 2.49465e-11, 2.485632e-11, 2.492689e-11, 2.479838e-11, 
    2.487027e-11, 2.491162e-11, 2.507144e-11, 2.510663e-11, 2.513923e-11, 
    2.520367e-11, 2.528643e-11, 2.543177e-11, 2.555844e-11, 2.567425e-11, 
    2.566576e-11, 2.566875e-11, 2.569462e-11, 2.563053e-11, 2.570515e-11, 
    2.571766e-11, 2.568492e-11, 2.587517e-11, 2.582078e-11, 2.587644e-11, 
    2.584103e-11, 2.495495e-11, 2.499867e-11, 2.497504e-11, 2.501948e-11, 
    2.498816e-11, 2.512746e-11, 2.516927e-11, 2.536521e-11, 2.528479e-11, 
    2.541286e-11, 2.52978e-11, 2.531817e-11, 2.541698e-11, 2.530403e-11, 
    2.555142e-11, 2.538357e-11, 2.569562e-11, 2.552768e-11, 2.570615e-11, 
    2.567375e-11, 2.572743e-11, 2.577551e-11, 2.583606e-11, 2.594784e-11, 
    2.592196e-11, 2.601554e-11, 2.506391e-11, 2.512069e-11, 2.511572e-11, 
    2.517519e-11, 2.521919e-11, 2.531467e-11, 2.546797e-11, 2.541031e-11, 
    2.551624e-11, 2.553751e-11, 2.53766e-11, 2.547533e-11, 2.515873e-11, 
    2.520977e-11, 2.51794e-11, 2.506837e-11, 2.542355e-11, 2.524108e-11, 
    2.557833e-11, 2.547928e-11, 2.576865e-11, 2.56246e-11, 2.59077e-11, 
    2.602889e-11, 2.614323e-11, 2.627683e-11, 2.515172e-11, 2.511312e-11, 
    2.518227e-11, 2.527797e-11, 2.536695e-11, 2.548531e-11, 2.549745e-11, 
    2.551963e-11, 2.557716e-11, 2.562554e-11, 2.552662e-11, 2.563768e-11, 
    2.522155e-11, 2.543942e-11, 2.509851e-11, 2.520099e-11, 2.527234e-11, 
    2.524106e-11, 2.540373e-11, 2.544209e-11, 2.559815e-11, 2.551746e-11, 
    2.599894e-11, 2.578562e-11, 2.637879e-11, 2.621266e-11, 2.509963e-11, 
    2.51516e-11, 2.533265e-11, 2.524647e-11, 2.549324e-11, 2.555406e-11, 
    2.560357e-11, 2.566683e-11, 2.567369e-11, 2.57112e-11, 2.564973e-11, 
    2.570878e-11, 2.548557e-11, 2.558526e-11, 2.531198e-11, 2.53784e-11, 
    2.534785e-11, 2.531432e-11, 2.541783e-11, 2.552817e-11, 2.553058e-11, 
    2.556598e-11, 2.566571e-11, 2.549424e-11, 2.602641e-11, 2.569732e-11, 
    2.52083e-11, 2.530848e-11, 2.532285e-11, 2.528402e-11, 2.554796e-11, 
    2.545223e-11, 2.571029e-11, 2.564049e-11, 2.57549e-11, 2.569803e-11, 
    2.568966e-11, 2.561668e-11, 2.557126e-11, 2.545661e-11, 2.536344e-11, 
    2.528966e-11, 2.530681e-11, 2.538789e-11, 2.553493e-11, 2.567429e-11, 
    2.564374e-11, 2.57462e-11, 2.547532e-11, 2.558879e-11, 2.55449e-11, 
    2.565938e-11, 2.540876e-11, 2.562199e-11, 2.535432e-11, 2.537777e-11, 
    2.545034e-11, 2.559645e-11, 2.562889e-11, 2.566343e-11, 2.564213e-11, 
    2.553868e-11, 2.552176e-11, 2.544858e-11, 2.542836e-11, 2.537267e-11, 
    2.532656e-11, 2.536867e-11, 2.541291e-11, 2.553874e-11, 2.565226e-11, 
    2.577619e-11, 2.580656e-11, 2.595147e-11, 2.583342e-11, 2.602823e-11, 
    2.586248e-11, 2.614964e-11, 2.563443e-11, 2.585771e-11, 2.545366e-11, 
    2.549711e-11, 2.557572e-11, 2.575635e-11, 2.565885e-11, 2.577292e-11, 
    2.55211e-11, 2.539066e-11, 2.5357e-11, 2.529413e-11, 2.535844e-11, 
    2.535321e-11, 2.541478e-11, 2.539499e-11, 2.554292e-11, 2.546344e-11, 
    2.568943e-11, 2.577203e-11, 2.600571e-11, 2.61492e-11, 2.629555e-11, 
    2.63602e-11, 2.637989e-11, 2.638812e-11,
  2.659464e-11, 2.673652e-11, 2.670893e-11, 2.682349e-11, 2.675994e-11, 
    2.683497e-11, 2.66234e-11, 2.674214e-11, 2.666633e-11, 2.660742e-11, 
    2.704622e-11, 2.682861e-11, 2.727304e-11, 2.713378e-11, 2.748409e-11, 
    2.725134e-11, 2.753111e-11, 2.747742e-11, 2.763924e-11, 2.759285e-11, 
    2.780007e-11, 2.766066e-11, 2.790775e-11, 2.776678e-11, 2.77888e-11, 
    2.765606e-11, 2.68724e-11, 2.701909e-11, 2.686371e-11, 2.688461e-11, 
    2.687523e-11, 2.676124e-11, 2.670382e-11, 2.658383e-11, 2.660561e-11, 
    2.669376e-11, 2.689401e-11, 2.6826e-11, 2.699758e-11, 2.69937e-11, 
    2.71851e-11, 2.709875e-11, 2.742112e-11, 2.732939e-11, 2.759479e-11, 
    2.752796e-11, 2.759164e-11, 2.757233e-11, 2.759189e-11, 2.74939e-11, 
    2.753587e-11, 2.744971e-11, 2.71149e-11, 2.721315e-11, 2.692045e-11, 
    2.67449e-11, 2.66286e-11, 2.654614e-11, 2.655779e-11, 2.658e-11, 
    2.669428e-11, 2.680189e-11, 2.688399e-11, 2.693895e-11, 2.699314e-11, 
    2.715729e-11, 2.724439e-11, 2.743967e-11, 2.740443e-11, 2.746416e-11, 
    2.752132e-11, 2.761731e-11, 2.760151e-11, 2.764382e-11, 2.746261e-11, 
    2.758298e-11, 2.738435e-11, 2.743863e-11, 2.700775e-11, 2.684435e-11, 
    2.677488e-11, 2.671423e-11, 2.656675e-11, 2.666856e-11, 2.662841e-11, 
    2.672399e-11, 2.678477e-11, 2.675471e-11, 2.694046e-11, 2.686819e-11, 
    2.724955e-11, 2.708507e-11, 2.751465e-11, 2.741166e-11, 2.753935e-11, 
    2.747418e-11, 2.758587e-11, 2.748534e-11, 2.765958e-11, 2.769755e-11, 
    2.76716e-11, 2.777138e-11, 2.747977e-11, 2.759163e-11, 2.675386e-11, 
    2.675876e-11, 2.678161e-11, 2.668121e-11, 2.667508e-11, 2.658323e-11, 
    2.666497e-11, 2.669979e-11, 2.67883e-11, 2.684068e-11, 2.689052e-11, 
    2.700019e-11, 2.712282e-11, 2.729465e-11, 2.741833e-11, 2.750133e-11, 
    2.745044e-11, 2.749537e-11, 2.744514e-11, 2.742161e-11, 2.768331e-11, 
    2.753625e-11, 2.775702e-11, 2.774479e-11, 2.764482e-11, 2.774617e-11, 
    2.676221e-11, 2.6734e-11, 2.663612e-11, 2.671271e-11, 2.657323e-11, 
    2.665126e-11, 2.669615e-11, 2.686967e-11, 2.690787e-11, 2.694327e-11, 
    2.701327e-11, 2.710316e-11, 2.726109e-11, 2.739876e-11, 2.752465e-11, 
    2.751542e-11, 2.751867e-11, 2.75468e-11, 2.747711e-11, 2.755824e-11, 
    2.757186e-11, 2.753625e-11, 2.774315e-11, 2.7684e-11, 2.774453e-11, 
    2.770601e-11, 2.674317e-11, 2.679065e-11, 2.676499e-11, 2.681324e-11, 
    2.677923e-11, 2.693051e-11, 2.697592e-11, 2.718877e-11, 2.710139e-11, 
    2.724054e-11, 2.711552e-11, 2.713765e-11, 2.724503e-11, 2.712228e-11, 
    2.739113e-11, 2.720872e-11, 2.754789e-11, 2.736534e-11, 2.755934e-11, 
    2.75241e-11, 2.758247e-11, 2.763476e-11, 2.770062e-11, 2.782222e-11, 
    2.779405e-11, 2.789587e-11, 2.686149e-11, 2.692314e-11, 2.691774e-11, 
    2.698233e-11, 2.703012e-11, 2.713384e-11, 2.730043e-11, 2.723775e-11, 
    2.735288e-11, 2.7376e-11, 2.720113e-11, 2.730843e-11, 2.696445e-11, 
    2.701991e-11, 2.69869e-11, 2.686633e-11, 2.725216e-11, 2.705391e-11, 
    2.742037e-11, 2.731271e-11, 2.76273e-11, 2.747068e-11, 2.777855e-11, 
    2.791041e-11, 2.803482e-11, 2.818029e-11, 2.695684e-11, 2.691492e-11, 
    2.699002e-11, 2.709399e-11, 2.719064e-11, 2.731927e-11, 2.733246e-11, 
    2.735657e-11, 2.74191e-11, 2.747169e-11, 2.736417e-11, 2.748488e-11, 
    2.703272e-11, 2.72694e-11, 2.689906e-11, 2.701036e-11, 2.708786e-11, 
    2.705389e-11, 2.72306e-11, 2.727229e-11, 2.744193e-11, 2.735421e-11, 
    2.787783e-11, 2.764577e-11, 2.829129e-11, 2.811041e-11, 2.690027e-11, 
    2.695671e-11, 2.715339e-11, 2.705976e-11, 2.732788e-11, 2.739399e-11, 
    2.74478e-11, 2.751659e-11, 2.752404e-11, 2.756483e-11, 2.7498e-11, 
    2.75622e-11, 2.731954e-11, 2.74279e-11, 2.713091e-11, 2.720309e-11, 
    2.716988e-11, 2.713346e-11, 2.724593e-11, 2.736586e-11, 2.736846e-11, 
    2.740695e-11, 2.751542e-11, 2.732897e-11, 2.790774e-11, 2.754978e-11, 
    2.701829e-11, 2.712713e-11, 2.714273e-11, 2.710054e-11, 2.738736e-11, 
    2.728332e-11, 2.756384e-11, 2.748794e-11, 2.761234e-11, 2.75505e-11, 
    2.75414e-11, 2.746206e-11, 2.741268e-11, 2.728808e-11, 2.718684e-11, 
    2.710667e-11, 2.71253e-11, 2.72134e-11, 2.737321e-11, 2.752469e-11, 
    2.749148e-11, 2.760288e-11, 2.730841e-11, 2.743174e-11, 2.738404e-11, 
    2.750849e-11, 2.723608e-11, 2.746787e-11, 2.717692e-11, 2.72024e-11, 
    2.728126e-11, 2.744008e-11, 2.747533e-11, 2.75129e-11, 2.748972e-11, 
    2.737728e-11, 2.735889e-11, 2.727935e-11, 2.725738e-11, 2.719685e-11, 
    2.714675e-11, 2.719252e-11, 2.724059e-11, 2.737734e-11, 2.750074e-11, 
    2.76355e-11, 2.766853e-11, 2.782619e-11, 2.769777e-11, 2.790973e-11, 
    2.772941e-11, 2.804184e-11, 2.748139e-11, 2.772419e-11, 2.728486e-11, 
    2.733209e-11, 2.741755e-11, 2.761394e-11, 2.75079e-11, 2.763195e-11, 
    2.735817e-11, 2.721642e-11, 2.717983e-11, 2.711153e-11, 2.718139e-11, 
    2.717571e-11, 2.724261e-11, 2.722111e-11, 2.738189e-11, 2.729549e-11, 
    2.754117e-11, 2.763098e-11, 2.788518e-11, 2.804134e-11, 2.820064e-11, 
    2.827104e-11, 2.829248e-11, 2.830144e-11,
  2.832222e-11, 2.847651e-11, 2.84465e-11, 2.857113e-11, 2.850197e-11, 
    2.858361e-11, 2.835348e-11, 2.848263e-11, 2.840016e-11, 2.833611e-11, 
    2.881361e-11, 2.85767e-11, 2.906068e-11, 2.890893e-11, 2.929079e-11, 
    2.903703e-11, 2.934207e-11, 2.928348e-11, 2.946003e-11, 2.940941e-11, 
    2.963566e-11, 2.948341e-11, 2.975325e-11, 2.959928e-11, 2.962334e-11, 
    2.947839e-11, 2.862433e-11, 2.878407e-11, 2.861487e-11, 2.863763e-11, 
    2.862742e-11, 2.850339e-11, 2.844095e-11, 2.831046e-11, 2.833413e-11, 
    2.843e-11, 2.864786e-11, 2.857385e-11, 2.876059e-11, 2.875637e-11, 
    2.896483e-11, 2.887076e-11, 2.922209e-11, 2.912206e-11, 2.941152e-11, 
    2.933861e-11, 2.940809e-11, 2.938702e-11, 2.940837e-11, 2.930147e-11, 
    2.934725e-11, 2.925326e-11, 2.888836e-11, 2.899539e-11, 2.867664e-11, 
    2.848564e-11, 2.835913e-11, 2.826949e-11, 2.828216e-11, 2.83063e-11, 
    2.843056e-11, 2.854761e-11, 2.863695e-11, 2.869676e-11, 2.875576e-11, 
    2.893456e-11, 2.902945e-11, 2.924232e-11, 2.920388e-11, 2.926903e-11, 
    2.933136e-11, 2.94361e-11, 2.941886e-11, 2.946503e-11, 2.926733e-11, 
    2.939866e-11, 2.918199e-11, 2.924118e-11, 2.877172e-11, 2.859381e-11, 
    2.851826e-11, 2.845226e-11, 2.82919e-11, 2.840259e-11, 2.835893e-11, 
    2.846287e-11, 2.852898e-11, 2.849628e-11, 2.86984e-11, 2.861975e-11, 
    2.903507e-11, 2.885588e-11, 2.932409e-11, 2.921177e-11, 2.935104e-11, 
    2.927995e-11, 2.94018e-11, 2.929212e-11, 2.948224e-11, 2.952369e-11, 
    2.949536e-11, 2.960428e-11, 2.928605e-11, 2.940808e-11, 2.849536e-11, 
    2.850069e-11, 2.852555e-11, 2.841635e-11, 2.840968e-11, 2.83098e-11, 
    2.839868e-11, 2.843655e-11, 2.853283e-11, 2.858982e-11, 2.864405e-11, 
    2.876343e-11, 2.8897e-11, 2.908422e-11, 2.921904e-11, 2.930956e-11, 
    2.925405e-11, 2.930306e-11, 2.924827e-11, 2.922261e-11, 2.950815e-11, 
    2.934767e-11, 2.958861e-11, 2.957526e-11, 2.946613e-11, 2.957676e-11, 
    2.850444e-11, 2.847376e-11, 2.836731e-11, 2.84506e-11, 2.829894e-11, 
    2.838378e-11, 2.843261e-11, 2.862137e-11, 2.866294e-11, 2.870147e-11, 
    2.877767e-11, 2.887557e-11, 2.904764e-11, 2.91977e-11, 2.9335e-11, 
    2.932493e-11, 2.932847e-11, 2.935916e-11, 2.928315e-11, 2.937165e-11, 
    2.938651e-11, 2.934766e-11, 2.957347e-11, 2.950889e-11, 2.957497e-11, 
    2.953292e-11, 2.848373e-11, 2.853538e-11, 2.850746e-11, 2.855996e-11, 
    2.852297e-11, 2.868759e-11, 2.873703e-11, 2.896884e-11, 2.887364e-11, 
    2.902525e-11, 2.888903e-11, 2.891314e-11, 2.903017e-11, 2.889639e-11, 
    2.918941e-11, 2.899059e-11, 2.936035e-11, 2.91613e-11, 2.937285e-11, 
    2.93344e-11, 2.939808e-11, 2.945515e-11, 2.952703e-11, 2.965982e-11, 
    2.962906e-11, 2.974026e-11, 2.861245e-11, 2.867957e-11, 2.867367e-11, 
    2.874398e-11, 2.879603e-11, 2.890898e-11, 2.90905e-11, 2.90222e-11, 
    2.914767e-11, 2.917288e-11, 2.898228e-11, 2.909923e-11, 2.872453e-11, 
    2.878492e-11, 2.874897e-11, 2.861774e-11, 2.903791e-11, 2.882195e-11, 
    2.922127e-11, 2.910389e-11, 2.944701e-11, 2.927615e-11, 2.961212e-11, 
    2.975618e-11, 2.989211e-11, 3.005119e-11, 2.871624e-11, 2.867061e-11, 
    2.875235e-11, 2.886559e-11, 2.897087e-11, 2.911104e-11, 2.912541e-11, 
    2.915171e-11, 2.921988e-11, 2.927724e-11, 2.916e-11, 2.929162e-11, 
    2.87989e-11, 2.905669e-11, 2.865335e-11, 2.877453e-11, 2.885892e-11, 
    2.88219e-11, 2.90144e-11, 2.905983e-11, 2.924478e-11, 2.914912e-11, 
    2.972058e-11, 2.946719e-11, 3.01726e-11, 2.997477e-11, 2.865466e-11, 
    2.871609e-11, 2.893029e-11, 2.882829e-11, 2.912042e-11, 2.919251e-11, 
    2.925117e-11, 2.932622e-11, 2.933434e-11, 2.937884e-11, 2.930592e-11, 
    2.937596e-11, 2.911135e-11, 2.922948e-11, 2.890579e-11, 2.898443e-11, 
    2.894824e-11, 2.890857e-11, 2.90311e-11, 2.916184e-11, 2.916467e-11, 
    2.920664e-11, 2.9325e-11, 2.912161e-11, 2.975331e-11, 2.936249e-11, 
    2.878314e-11, 2.890169e-11, 2.891867e-11, 2.887271e-11, 2.918528e-11, 
    2.907186e-11, 2.937776e-11, 2.929496e-11, 2.943068e-11, 2.936321e-11, 
    2.935328e-11, 2.926673e-11, 2.921289e-11, 2.907705e-11, 2.896672e-11, 
    2.887938e-11, 2.889968e-11, 2.899566e-11, 2.916986e-11, 2.933506e-11, 
    2.929883e-11, 2.942036e-11, 2.90992e-11, 2.923368e-11, 2.918166e-11, 
    2.931737e-11, 2.902038e-11, 2.927313e-11, 2.89559e-11, 2.898367e-11, 
    2.906961e-11, 2.924279e-11, 2.92812e-11, 2.932219e-11, 2.92969e-11, 
    2.917429e-11, 2.915423e-11, 2.906752e-11, 2.904359e-11, 2.897762e-11, 
    2.892304e-11, 2.89729e-11, 2.90253e-11, 2.917435e-11, 2.930893e-11, 
    2.945596e-11, 2.9492e-11, 2.966419e-11, 2.952396e-11, 2.975549e-11, 
    2.955855e-11, 2.989983e-11, 2.928785e-11, 2.95528e-11, 2.907353e-11, 
    2.912501e-11, 2.92182e-11, 2.943245e-11, 2.931674e-11, 2.94521e-11, 
    2.915345e-11, 2.899897e-11, 2.895908e-11, 2.888468e-11, 2.896078e-11, 
    2.895459e-11, 2.902749e-11, 2.900405e-11, 2.91793e-11, 2.908512e-11, 
    2.935303e-11, 2.945104e-11, 2.972859e-11, 2.989925e-11, 3.007342e-11, 
    3.015044e-11, 3.017389e-11, 3.01837e-11,
  2.87211e-11, 2.888357e-11, 2.885195e-11, 2.898328e-11, 2.891039e-11, 
    2.899644e-11, 2.8754e-11, 2.889002e-11, 2.880315e-11, 2.873571e-11, 
    2.923913e-11, 2.898915e-11, 2.950011e-11, 2.933973e-11, 2.974359e-11, 
    2.947512e-11, 2.979789e-11, 2.973583e-11, 2.992287e-11, 2.986921e-11, 
    3.010918e-11, 2.994765e-11, 3.023401e-11, 3.007056e-11, 3.009609e-11, 
    2.994233e-11, 2.903936e-11, 2.920793e-11, 2.902939e-11, 2.905339e-11, 
    2.904262e-11, 2.891189e-11, 2.884613e-11, 2.870871e-11, 2.873363e-11, 
    2.883458e-11, 2.906419e-11, 2.898613e-11, 2.918309e-11, 2.917863e-11, 
    2.939878e-11, 2.92994e-11, 2.967084e-11, 2.9565e-11, 2.987145e-11, 
    2.979421e-11, 2.986782e-11, 2.984549e-11, 2.986811e-11, 2.975488e-11, 
    2.980336e-11, 2.970383e-11, 2.9318e-11, 2.943109e-11, 2.909453e-11, 
    2.889322e-11, 2.875995e-11, 2.86656e-11, 2.867893e-11, 2.870435e-11, 
    2.883517e-11, 2.895848e-11, 2.905266e-11, 2.911575e-11, 2.917799e-11, 
    2.936685e-11, 2.94671e-11, 2.969227e-11, 2.965156e-11, 2.972054e-11, 
    2.978653e-11, 2.989751e-11, 2.987923e-11, 2.992818e-11, 2.971873e-11, 
    2.985783e-11, 2.962839e-11, 2.969104e-11, 2.919491e-11, 2.900718e-11, 
    2.892758e-11, 2.885802e-11, 2.868918e-11, 2.880571e-11, 2.875974e-11, 
    2.886918e-11, 2.893885e-11, 2.890438e-11, 2.911747e-11, 2.903452e-11, 
    2.947304e-11, 2.92837e-11, 2.977883e-11, 2.965992e-11, 2.980738e-11, 
    2.973208e-11, 2.986116e-11, 2.974497e-11, 2.994641e-11, 2.999038e-11, 
    2.996033e-11, 3.007586e-11, 2.973854e-11, 2.986782e-11, 2.890342e-11, 
    2.890904e-11, 2.893522e-11, 2.882021e-11, 2.881318e-11, 2.870802e-11, 
    2.880158e-11, 2.884147e-11, 2.894289e-11, 2.900297e-11, 2.906015e-11, 
    2.91861e-11, 2.932713e-11, 2.952499e-11, 2.966762e-11, 2.976344e-11, 
    2.970466e-11, 2.975655e-11, 2.969855e-11, 2.967138e-11, 2.99739e-11, 
    2.980382e-11, 3.005923e-11, 3.004506e-11, 2.992935e-11, 3.004665e-11, 
    2.891298e-11, 2.888065e-11, 2.876856e-11, 2.885626e-11, 2.869658e-11, 
    2.87859e-11, 2.883733e-11, 2.903625e-11, 2.908007e-11, 2.912072e-11, 
    2.920112e-11, 2.930448e-11, 2.948631e-11, 2.964504e-11, 2.979038e-11, 
    2.977971e-11, 2.978347e-11, 2.981598e-11, 2.973547e-11, 2.982921e-11, 
    2.984496e-11, 2.980379e-11, 3.004316e-11, 2.997467e-11, 3.004476e-11, 
    3.000015e-11, 2.889116e-11, 2.894558e-11, 2.891617e-11, 2.89715e-11, 
    2.893251e-11, 2.91061e-11, 2.915826e-11, 2.940304e-11, 2.930245e-11, 
    2.946264e-11, 2.93187e-11, 2.934417e-11, 2.946788e-11, 2.932646e-11, 
    2.963627e-11, 2.942603e-11, 2.981724e-11, 2.960655e-11, 2.983048e-11, 
    2.978975e-11, 2.985721e-11, 2.99177e-11, 2.999391e-11, 3.013481e-11, 
    3.010215e-11, 3.02202e-11, 2.902683e-11, 2.909762e-11, 2.909139e-11, 
    2.916557e-11, 2.92205e-11, 2.933976e-11, 2.953163e-11, 2.94594e-11, 
    2.959209e-11, 2.961877e-11, 2.941721e-11, 2.954087e-11, 2.914506e-11, 
    2.92088e-11, 2.917084e-11, 2.903241e-11, 2.947603e-11, 2.924789e-11, 
    2.966997e-11, 2.954579e-11, 2.990907e-11, 2.972808e-11, 3.008418e-11, 
    3.023715e-11, 3.038154e-11, 3.055078e-11, 2.91363e-11, 2.908815e-11, 
    2.91744e-11, 2.929396e-11, 2.940516e-11, 2.955335e-11, 2.956854e-11, 
    2.959636e-11, 2.966849e-11, 2.972921e-11, 2.960516e-11, 2.974444e-11, 
    2.922359e-11, 2.949588e-11, 2.906996e-11, 2.919784e-11, 2.928691e-11, 
    2.924782e-11, 2.945115e-11, 2.949919e-11, 2.969487e-11, 2.959362e-11, 
    3.019935e-11, 2.993049e-11, 3.068002e-11, 3.046947e-11, 2.907134e-11, 
    2.913614e-11, 2.936229e-11, 2.925456e-11, 2.956326e-11, 2.963953e-11, 
    2.970162e-11, 2.978109e-11, 2.978968e-11, 2.983683e-11, 2.975959e-11, 
    2.983378e-11, 2.955367e-11, 2.967866e-11, 2.933639e-11, 2.941949e-11, 
    2.938124e-11, 2.933933e-11, 2.946881e-11, 2.96071e-11, 2.961007e-11, 
    2.965449e-11, 2.977988e-11, 2.956452e-11, 3.023414e-11, 2.981957e-11, 
    2.920689e-11, 2.93321e-11, 2.935001e-11, 2.930145e-11, 2.963188e-11, 
    2.951191e-11, 2.983568e-11, 2.974798e-11, 2.989176e-11, 2.982026e-11, 
    2.980975e-11, 2.971809e-11, 2.96611e-11, 2.95174e-11, 2.940078e-11, 
    2.93085e-11, 2.932994e-11, 2.943137e-11, 2.961558e-11, 2.979045e-11, 
    2.97521e-11, 2.988082e-11, 2.954082e-11, 2.968311e-11, 2.962807e-11, 
    2.977172e-11, 2.945748e-11, 2.972493e-11, 2.938934e-11, 2.941868e-11, 
    2.950953e-11, 2.969277e-11, 2.973341e-11, 2.977682e-11, 2.975003e-11, 
    2.962026e-11, 2.959904e-11, 2.950732e-11, 2.948202e-11, 2.941229e-11, 
    2.935462e-11, 2.94073e-11, 2.946269e-11, 2.962032e-11, 2.976279e-11, 
    2.991856e-11, 2.995676e-11, 3.013948e-11, 2.999068e-11, 3.023646e-11, 
    3.002743e-11, 3.038982e-11, 2.974049e-11, 3.002129e-11, 2.951367e-11, 
    2.956812e-11, 2.966674e-11, 2.989367e-11, 2.977104e-11, 2.991448e-11, 
    2.95982e-11, 2.943487e-11, 2.939269e-11, 2.93141e-11, 2.939449e-11, 
    2.938795e-11, 2.946499e-11, 2.944022e-11, 2.962556e-11, 2.952592e-11, 
    2.980948e-11, 2.991335e-11, 3.020782e-11, 3.038916e-11, 3.057441e-11, 
    3.065641e-11, 3.068139e-11, 3.069184e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
